// -----------------------------------------------------------------------------
//Actel Corporation Proprietary and Confidential
//Copyright 2008 Actel Corporation. All rights reserved.
//
//ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
//ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
//IN ADVANCE IN WRITING.
//
//Description:  CoreFFT RTL 
//              Customized Twiddle Coefficients 
//
//Revision Information:
//Date         Description
//05Nov2009    Initial Release 
//
//SVN Revision Information:
//SVN $Revision: $
//SVN $Data: $
//
//Resolved SARs
//SAR     Date    Who         Description
//
//Notes:

`timescale 1 ns/100 ps

module COREFFT_C0_COREFFT_C0_0_twiddle (A,T);
  parameter TDWIDTH = 16;
  parameter LOGPTS  = 5;

  input	[LOGPTS-2:0]	A;	// Address
  output reg [TDWIDTH-1:0]	T;	// Table output

  always @ (A)
    case (A) // synopsys parallel_case
      11'h0: T=64'b0000000000000000000000000000000001111111111111111111111111111111;  //     0 2147483647
      11'h1: T=64'b1111111111001101101111000000101101111111111111111111011000100000;  // -3294197 2147481120
      11'h2: T=64'b1111111110011011011110000001110101111111111111111101100010000101;  // -6588387 2147473541
      11'h3: T=64'b1111111101101001001101000011111101111111111111111010011100101011;  // -9882561 2147460907
      11'h4: T=64'b1111111100110110111100000111100001111111111111110110001000010101;  // -13176712 2147443221
      11'h5: T=64'b1111111100000100101011001101000001111111111111110000100101000010;  // -16470832 2147420482
      11'h6: T=64'b1111111011010010011010010100111101111111111111101001110010110001;  // -19764913 2147392689
      11'h7: T=64'b1111111010100000001001011111110101111111111111100001110001100100;  // -23058947 2147359844
      11'h8: T=64'b1111111001101101111000101110000001111111111111011000100001011001;  // -26352928 2147321945
      11'h9: T=64'b1111111000111011101000000000001001111111111111001110000010010010;  // -29646846 2147278994
      11'ha: T=64'b1111111000001001010111010110100101111111111111000010010100001110;  // -32940695 2147230990
      11'hb: T=64'b1111110111010111000110110001111001111111111110110101010111001101;  // -36234466 2147177933
      11'hc: T=64'b1111110110100100110110010010100101111111111110100111001011010000;  // -39528151 2147119824
      11'hd: T=64'b1111110101110010100101111001000001111111111110010111110000010111;  // -42821744 2147056663
      11'he: T=64'b1111110101000000010101100101110001111111111110000111000110100001;  // -46115236 2146988449
      11'hf: T=64'b1111110100001110000101011001010001111111111101110101001101101111;  // -49408620 2146915183
      11'h10: T=64'b1111110011011011110101010100000101111111111101100010000110000001;  // -52701887 2146836865
      11'h11: T=64'b1111110010101001100101010110101001111111111101001101101111011000;  // -55995030 2146753496
      11'h12: T=64'b1111110001110111010101100001011001111111111100111000001001110011;  // -59288042 2146665075
      11'h13: T=64'b1111110001000101000101110100111001111111111100100001010101010010;  // -62580914 2146571602
      11'h14: T=64'b1111110000010010110110010001101001111111111100001001010001110111;  // -65873638 2146473079
      11'h15: T=64'b1111101111100000100110111000000001111111111011101111111111100000;  // -69166208 2146369504
      11'h16: T=64'b1111101110101110010111101000100101111111111011010101011110010000;  // -72458615 2146260880
      11'h17: T=64'b1111101101111100001000100011110101111111111010111001101110000100;  // -75750851 2146147204
      11'h18: T=64'b1111101101001001111001101010001101111111111010011100101110111111;  // -79042909 2146028479
      11'h19: T=64'b1111101100010111101010111100001001111111111001111110100001000000;  // -82334782 2145904704
      11'h1a: T=64'b1111101011100101011100011010010001111111111001011111000100000111;  // -85626460 2145775879
      11'h1b: T=64'b1111101010110011001110000100111101111111111000111110011000010101;  // -88917937 2145642005
      11'h1c: T=64'b1111101010000000111111111100101101111111111000011100011101101010;  // -92209205 2145503082
      11'h1d: T=64'b1111101001001110110010000010000101111111110111111001010100000111;  // -95500255 2145359111
      11'h1e: T=64'b1111101000011100100100010101011101111111110111010100111011101011;  // -98791081 2145210091
      11'h1f: T=64'b1111100111101010010110110111010101111111110110101111010100011000;  // -102081675 2145056024
      11'h20: T=64'b1111100110111000001001101000010001111111110110001000011110001101;  // -105372028 2144896909
      11'h21: T=64'b1111100110000101111100101000101001111111110101100000011001001011;  // -108662134 2144732747
      11'h22: T=64'b1111100101010011101111111001000101111111110100110111000101010010;  // -111951983 2144563538
      11'h23: T=64'b1111100100100001100011011001111001111111110100001100100010100010;  // -115241570 2144389282
      11'h24: T=64'b1111100011101111010111001011101101111111110011100000110000111101;  // -118530885 2144209981
      11'h25: T=64'b1111100010111101001011001110111101111111110010110011110000100010;  // -121819921 2144025634
      11'h26: T=64'b1111100010001010111111100100001001111111110010000101100001010011;  // -125108670 2143836243
      11'h27: T=64'b1111100001011000110100001011101101111111110001010110000011001110;  // -128397125 2143641806
      11'h28: T=64'b1111100000100110101001000110001001111111110000100101010110010101;  // -131685278 2143442325
      11'h29: T=64'b1111011111110100011110010011111001111111101111110011011010101001;  // -134973122 2143237801
      11'h2a: T=64'b1111011111000010010011110101100101111111101111000000010000001001;  // -138260647 2143028233
      11'h2b: T=64'b1111011110010000001001101011100101111111101110001011110110110111;  // -141547847 2142813623
      11'h2c: T=64'b1111011101011101111111110110011001111111101101010110001110110010;  // -144834714 2142593970
      11'h2d: T=64'b1111011100101011110110010110011101111111101100011111010111111011;  // -148121241 2142369275
      11'h2e: T=64'b1111011011111001101101001100011001111111101011100111010010010100;  // -151407418 2142139540
      11'h2f: T=64'b1111011011000111100100011000100001111111101010101101111101111011;  // -154693240 2141904763
      11'h30: T=64'b1111011010010101011011111011011101111111101001110011011010110011;  // -157978697 2141664947
      11'h31: T=64'b1111011001100011010011110101100101111111101000110111101000111011;  // -161263783 2141420091
      11'h32: T=64'b1111011000110001001100000111011101111111100111111010101000010100;  // -164548489 2141170196
      11'h33: T=64'b1111010111111111000100110001100001111111100110111100011000111111;  // -167832808 2140915263
      11'h34: T=64'b1111010111001100111101110100010001111111100101111100111010111100;  // -171116732 2140655292
      11'h35: T=64'b1111010110011010110111010000001001111111100100111100001110001011;  // -174400254 2140390283
      11'h36: T=64'b1111010101101000110001000101101101111111100011111010010010101111;  // -177683365 2140120239
      11'h37: T=64'b1111010100110110101011010101011001111111100010110111001000100110;  // -180966058 2139845158
      11'h38: T=64'b1111010100000100100101111111101101111111100001110010101111110010;  // -184248325 2139565042
      11'h39: T=64'b1111010011010010100001000101000101111111100000101101001000010011;  // -187530159 2139279891
      11'h3a: T=64'b1111010010100000011100100110000101111111011111100110010010001011;  // -190811551 2138989707
      11'h3b: T=64'b1111010001101110011000100011001001111111011110011110001101011001;  // -194092494 2138694489
      11'h3c: T=64'b1111010000111100010100111100101101111111011101010100111001111111;  // -197372981 2138394239
      11'h3d: T=64'b1111010000001010010001110011010101111111011100001010010111111101;  // -200653003 2138088957
      11'h3e: T=64'b1111001111011000001111000111011101111111011010111110100111010011;  // -203932553 2137778643
      11'h3f: T=64'b1111001110100110001100111001100101111111011001110001101000000100;  // -207211623 2137463300
      11'h40: T=64'b1111001101110100001011001010001001111111011000100011011010001110;  // -210490206 2137142926
      11'h41: T=64'b1111001101000010001001111001101101111111010111010011111101110100;  // -213768293 2136817524
      11'h42: T=64'b1111001100010000001001001000101101111111010110000011010010110110;  // -217045877 2136487094
      11'h43: T=64'b1111001011011110001000110111100101111111010100110001011001010100;  // -220322951 2136151636
      11'h44: T=64'b1111001010101100001001000110111001111111010011011110010001010000;  // -223599506 2135811152
      11'h45: T=64'b1111001001111010001001110111000101111111010010001001111010101001;  // -226875535 2135465641
      11'h46: T=64'b1111001001001000001011001000101001111111010000110100010101100010;  // -230151030 2135115106
      11'h47: T=64'b1111001000010110001100111100000101111111001111011101100001111011;  // -233425983 2134759547
      11'h48: T=64'b1111000111100100001111010001110001111111001110000101011111110101;  // -236700388 2134398965
      11'h49: T=64'b1111000110110010010010001010010101111111001100101100001111010000;  // -239974235 2134033360
      11'h4a: T=64'b1111000110000000010101100110001101111111001011010001110000001101;  // -243247517 2133662733
      11'h4b: T=64'b1111000101001110011001100101110001111111001001110110000010101110;  // -246520228 2133287086
      11'h4c: T=64'b1111000100011100011110001001101001111111001000011001000110110011;  // -249792358 2132906419
      11'h4d: T=64'b1111000011101010100011010010010001111111000110111010111100011101;  // -253063900 2132520733
      11'h4e: T=64'b1111000010111000101001000000000101111111000101011011100011101101;  // -256334847 2132130029
      11'h4f: T=64'b1111000010000110101111010011101001111111000011111010111100100100;  // -259605190 2131734308
      11'h50: T=64'b1111000001010100110110001101010101111111000010011001000111000011;  // -262874923 2131333571
      11'h51: T=64'b1111000000100010111101101101101101111111000000110110000011001010;  // -266144037 2130927818
      11'h52: T=64'b1110111111110001000101110101001101111110111111010001110000111011;  // -269412525 2130517051
      11'h53: T=64'b1110111110111111001110100100010101111110111101101100010000010111;  // -272680379 2130101271
      11'h54: T=64'b1110111110001101010111111011100001111110111100000101100001011111;  // -275947592 2129680479
      11'h55: T=64'b1110111101011011100001111011010101111110111010011101100100010011;  // -279214155 2129254675
      11'h56: T=64'b1110111100101001101100100100001101111110111000110100011000110101;  // -282480061 2128823861
      11'h57: T=64'b1110111011110111110111110110101001111110110111001001111111000101;  // -285745302 2128388037
      11'h58: T=64'b1110111011000110000011110011000101111110110101011110010111000101;  // -289009871 2127947205
      11'h59: T=64'b1110111010010100010000011010000001111110110011110001100000110110;  // -292273760 2127501366
      11'h5a: T=64'b1110111001100010011101101011111101111110110010000011011100011001;  // -295536961 2127050521
      11'h5b: T=64'b1110111000110000101011101001011001111110110000010100001001101111;  // -298799466 2126594671
      11'h5c: T=64'b1110110111111110111010010010101101111110101110100011101000111000;  // -302061269 2126133816
      11'h5d: T=64'b1110110111001101001001101000011101111110101100110001111001110111;  // -305322361 2125667959
      11'h5e: T=64'b1110110110011011011001101011001001111110101010111110111100101011;  // -308582734 2125197099
      11'h5f: T=64'b1110110101101001101010011011001101111110101001001010110001010111;  // -311842381 2124721239
      11'h60: T=64'b1110110100110111111011111001001001111110100111010101010111111011;  // -315101294 2124240379
      11'h61: T=64'b1110110100000110001110000101011001111110100101011110110000011001;  // -318359466 2123754521
      11'h62: T=64'b1110110011010100100001000000011101111110100011100110111010110001;  // -321616889 2123263665
      11'h63: T=64'b1110110010100010110100101010110101111110100001101101110111000101;  // -324873555 2122767813
      11'h64: T=64'b1110110001110001001001000100111101111110011111110011100101010110;  // -328129457 2122266966
      11'h65: T=64'b1110110000111111011110001111011001111110011101111000000101100101;  // -331384586 2121761125
      11'h66: T=64'b1110110000001101110100001010100001111110011011111011010111110011;  // -334638936 2121250291
      11'h67: T=64'b1110101111011100001010110110111001111110011001111101011100000010;  // -337892498 2120734466
      11'h68: T=64'b1110101110101010100010010100111101111110010111111110010010010010;  // -341145265 2120213650
      11'h69: T=64'b1110101101111000111010100101001101111110010101111101111010100110;  // -344397229 2119687846
      11'h6a: T=64'b1110101101000111010011101000000101111110010011111100010100111101;  // -347648383 2119157053
      11'h6b: T=64'b1110101100010101101101011110000101111110010001111001100001011010;  // -350898719 2118621274
      11'h6c: T=64'b1110101011100100001000000111101101111110001111110101011111111110;  // -354148229 2118080510
      11'h6d: T=64'b1110101010110010100011100101011001111110001101110000010000101001;  // -357396906 2117534761
      11'h6e: T=64'b1110101010000000111111110111101001111110001011101001110011011110;  // -360644742 2116984030
      11'h6f: T=64'b1110101001001111011100111110111101111110001001100010001000011110;  // -363891729 2116428318
      11'h70: T=64'b1110101000011101111010111011110001111110000111011001001111101001;  // -367137860 2115867625
      11'h71: T=64'b1110100111101100011001101110100101111110000101001111001001000001;  // -370383127 2115301953
      11'h72: T=64'b1110100110111010111001010111110101111110000011000011110100101000;  // -373627523 2114731304
      11'h73: T=64'b1110100110001001011001111000000101111110000000110111010010011111;  // -376871039 2114155679
      11'h74: T=64'b1110100101010111111011001111101101111101111110101001100010100111;  // -380113669 2113575079
      11'h75: T=64'b1110100100100110011101011111010001111101111100011010100101000001;  // -383355404 2112989505
      11'h76: T=64'b1110100011110101000000100111001101111101111010001010011001101111;  // -386596237 2112398959
      11'h77: T=64'b1110100011000011100100101000000001111101110111111001000000110011;  // -389836160 2111803443
      11'h78: T=64'b1110100010010010001001100010001001111101110101100110011010001110;  // -393075166 2111202958
      11'h79: T=64'b1110100001100000101111010110000101111101110011010010100110000000;  // -396313247 2110597504
      11'h7a: T=64'b1110100000101111010110000100010001111101110000111101100100001100;  // -399550396 2109987084
      11'h7b: T=64'b1110011111111101111101101101010001111101101110100111010100110011;  // -402786604 2109371699
      11'h7c: T=64'b1110011111001100100110010001100001111101101100001111110111110111;  // -406021864 2108751351
      11'h7d: T=64'b1110011110011011001111110001011001111101101001110111001101011000;  // -409256170 2108126040
      11'h7e: T=64'b1110011101101001111010001101100001111101100111011101010101011001;  // -412489512 2107495769
      11'h7f: T=64'b1110011100111000100101100110010101111101100101000010001111111011;  // -415721883 2106860539
      11'h80: T=64'b1110011100000111010001111100010001111101100010100101111100111111;  // -418953276 2106220351
      11'h81: T=64'b1110011011010101111111001111110001111101100000001000011100100111;  // -422183684 2105575207
      11'h82: T=64'b1110011010100100101101100001011001111101011101101001101110110100;  // -425413098 2104925108
      11'h83: T=64'b1110011001110011011100110001101001111101011011001001110011101000;  // -428641510 2104270056
      11'h84: T=64'b1110011001000010001101000000110101111101011000101000101011000101;  // -431868915 2103610053
      11'h85: T=64'b1110011000010000111110001111100101111101010110000110010101001100;  // -435095303 2102945100
      11'h86: T=64'b1110010111011111110000011110010101111101010011100010110001111110;  // -438320667 2102275198
      11'h87: T=64'b1110010110101110100011101101100001111101010000111110000001011101;  // -441545000 2101600349
      11'h88: T=64'b1110010101111101010111111101101101111101001110011000000011101011;  // -444768293 2100920555
      11'h89: T=64'b1110010101001100001101001111001101111101001011110000111000101010;  // -447990541 2100235818
      11'h8a: T=64'b1110010100011011000011100010101001111101001001001000100000011010;  // -451211734 2099546138
      11'h8b: T=64'b1110010011101001111010111000011101111101000110011110111010111110;  // -454431865 2098851518
      11'h8c: T=64'b1110010010111000110011010001000101111101000011110100001000010111;  // -457650927 2098151959
      11'h8d: T=64'b1110010010000111101100101101000001111101000001001000001000100111;  // -460868912 2097447463
      11'h8e: T=64'b1110010001010110100111001100101101111100111110011010111011101111;  // -464085813 2096738031
      11'h8f: T=64'b1110010000100101100010110000101101111100111011101100100001110010;  // -467301621 2096023666
      11'h90: T=64'b1110001111110100011111011001011001111100111000111100111010110001;  // -470516330 2095304369
      11'h91: T=64'b1110001111000011011101000111010001111100110110001100000110101101;  // -473729932 2094580141
      11'h92: T=64'b1110001110010010011011111010110101111100110011011010000101101000;  // -476942419 2093850984
      11'h93: T=64'b1110001101100001011011110100100001111100110000100110110111100100;  // -480153784 2093116900
      11'h94: T=64'b1110001100110000011100110100110101111100101101110010011100100011;  // -483364019 2092377891
      11'h95: T=64'b1110001011111111011110111100010001111100101010111100110100100111;  // -486573116 2091633959
      11'h96: T=64'b1110001011001110100010001011001101111100101000000101111111110000;  // -489781069 2090885104
      11'h97: T=64'b1110001010011101100110100010001101111100100101001101111110000010;  // -492987869 2090131330
      11'h98: T=64'b1110001001101100101100000001101101111100100010010100101111011101;  // -496193509 2089372637
      11'h99: T=64'b1110001000111011110010101010001101111100011111011010010100000100;  // -499397981 2088609028
      11'h9a: T=64'b1110001000001010111010011100000101111100011100011110101011111000;  // -502601279 2087840504
      11'h9b: T=64'b1110000111011010000011010111111101111100011001100001110110111011;  // -505803393 2087067067
      11'h9c: T=64'b1110000110101001001101011110001001111100010110100011110101001111;  // -509004318 2086288719
      11'h9d: T=64'b1110000101111000011000101111001101111100010011100100100110110110;  // -512204045 2085505462
      11'h9e: T=64'b1110000101000111100101001011101001111100010000100100001011110001;  // -515402566 2084717297
      11'h9f: T=64'b1110000100010110110010110011110101111100001101100010100100000011;  // -518599875 2083924227
      11'ha0: T=64'b1110000011100110000001101000010101111100001010011111101111101101;  // -521795963 2083126253
      11'ha1: T=64'b1110000010110101010001101001100101111100000111011011101110110010;  // -524990823 2082323378
      11'ha2: T=64'b1110000010000100100010111000000001111100000100010110100001010010;  // -528184448 2081515602
      11'ha3: T=64'b1110000001010011110101010100000101111100000001010000000111010001;  // -531376831 2080702929
      11'ha4: T=64'b1110000000100011001000111110010101111011111110001000100000101111;  // -534567963 2079885359
      11'ha5: T=64'b1101111111110010011101110111001101111011111010111111101101101111;  // -537757837 2079062895
      11'ha6: T=64'b1101111111000001110011111111001101111011110111110101101110010011;  // -540946445 2078235539
      11'ha7: T=64'b1101111110010001001011010110101101111011110100101010100010011101;  // -544133781 2077403293
      11'ha8: T=64'b1101111101100000100011111110010001111011110001011110001010001111;  // -547319836 2076566159
      11'ha9: T=64'b1101111100101111111101110110010001111011101110010000100101101010;  // -550504604 2075724138
      11'haa: T=64'b1101111011111111011000111111010001111011101011000001110100110000;  // -553688076 2074877232
      11'hab: T=64'b1101111011001110110101011001101101111011100111110001110111100101;  // -556870245 2074025445
      11'hac: T=64'b1101111010011110010011000110000101111011100100100000101110001000;  // -560051103 2073168776
      11'had: T=64'b1101111001101101110010000100110001111011100001001110011000011110;  // -563230644 2072307230
      11'hae: T=64'b1101111000111101010010010110010001111011011101111010110110100111;  // -566408860 2071440807
      11'haf: T=64'b1101111000001100110011111011000101111011011010100110001000100110;  // -569585743 2070569510
      11'hb0: T=64'b1101110111011100010110110011101101111011010111010000001110011101;  // -572761285 2069693341
      11'hb1: T=64'b1101110110101011111011000000100001111011010011111001001000001101;  // -575935480 2068812301
      11'hb2: T=64'b1101110101111011100000100010000101111011010000100000110101111001;  // -579108319 2067926393
      11'hb3: T=64'b1101110101001011000111011000110001111011001101000111010111100100;  // -582279796 2067035620
      11'hb4: T=64'b1101110100011010101111100101000101111011001001101100101101001110;  // -585449903 2066139982
      11'hb5: T=64'b1101110011101010011001000111100001111011000110010000110110111011;  // -588618632 2065239483
      11'hb6: T=64'b1101110010111010000100000000100001111011000010110011110100101011;  // -591785976 2064334123
      11'hb7: T=64'b1101110010001001110000010000100101111010111111010101100110100011;  // -594951927 2063423907
      11'hb8: T=64'b1101110001011001011101111000001001111010111011110110001100100011;  // -598116478 2062508835
      11'hb9: T=64'b1101110000101001001100110111101001111010111000010101100110101101;  // -601279622 2061588909
      11'hba: T=64'b1101101111111000111101001111100101111010110100110011110101000100;  // -604441351 2060664132
      11'hbb: T=64'b1101101111001000101111000000011001111010110001010000110111101011;  // -607601658 2059734507
      11'hbc: T=64'b1101101110011000100010001010100101111010101101101100101110100011;  // -610760535 2058800035
      11'hbd: T=64'b1101101101101000010110101110100101111010101010000111011001101110;  // -613917975 2057860718
      11'hbe: T=64'b1101101100111000001100101100111001111010100110100000111001001111;  // -617073970 2056916559
      11'hbf: T=64'b1101101100001000000100000101111001111010100010111001001101000111;  // -620228514 2055967559
      11'hc0: T=64'b1101101011010111111100111010001101111010011111010000010101011010;  // -623381597 2055013722
      11'hc1: T=64'b1101101010100111110111001010001001111010011011100110010010001001;  // -626533214 2054055049
      11'hc2: T=64'b1101101001110111110010110110001101111010010111111011000011010111;  // -629683357 2053091543
      11'hc3: T=64'b1101101001000111101111111110111001111010010100001110101001000110;  // -632832018 2052123206
      11'hc4: T=64'b1101101000010111101110100100101001111010010000100001000011011000;  // -635979190 2051150040
      11'hc5: T=64'b1101100111100111101110100111111101111010001100110010010010001111;  // -639124865 2050172047
      11'hc6: T=64'b1101100110110111110000001001010001111010001001000010010101101110;  // -642269036 2049189230
      11'hc7: T=64'b1101100110000111110011001001000001111010000101010001001101110111;  // -645411696 2048201591
      11'hc8: T=64'b1101100101010111110111100111101101111010000001011110111010101100;  // -648552837 2047209132
      11'hc9: T=64'b1101100100100111111101100101101101111001111101101011011100010000;  // -651692453 2046211856
      11'hca: T=64'b1101100011111000000101000011101001111001111001110110110010100110;  // -654830534 2045209766
      11'hcb: T=64'b1101100011001000001110000001110101111001110110000000111101101110;  // -657967075 2044202862
      11'hcc: T=64'b1101100010011000011000100000110001111001110010001001111101101101;  // -661102068 2043191149
      11'hcd: T=64'b1101100001101000100100100000111101111001101110010001110010100011;  // -664235505 2042174627
      11'hce: T=64'b1101100000111000110010000010110101111001101010011000011100010101;  // -667367379 2041153301
      11'hcf: T=64'b1101100000001001000001000110111001111001100110011101111011000011;  // -670497682 2040127171
      11'hd0: T=64'b1101011111011001010001101101100001111001100010100010001110110000;  // -673626408 2039096240
      11'hd1: T=64'b1101011110101001100011110111001101111001011110100101010111100000;  // -676753549 2038060512
      11'hd2: T=64'b1101011101111001110111100100011101111001011010100111010101010011;  // -679879097 2037019987
      11'hd3: T=64'b1101011101001010001100110101101101111001010110101000001000001101;  // -683003045 2035974669
      11'hd4: T=64'b1101011100011010100011101011011001111001010010100111110000010001;  // -686125386 2034924561
      11'hd5: T=64'b1101011011101010111100000101111101111001001110100110001101100000;  // -689246113 2033869664
      11'hd6: T=64'b1101011010111011010110000101111001111001001010100011011111111101;  // -692365218 2032809981
      11'hd7: T=64'b1101011010001011110001101011101001111001000110011111100111101011;  // -695482694 2031745515
      11'hd8: T=64'b1101011001011100001110110111101101111001000010011010100100101100;  // -698598533 2030676268
      11'hd9: T=64'b1101011000101100101101101010100001111000111110010100010111000010;  // -701712728 2029602242
      11'hda: T=64'b1101010111111101001110000100100001111000111010001100111110110001;  // -704825272 2028523441
      11'hdb: T=64'b1101010111001101110000000110001101111000110110000100011011111010;  // -707936157 2027439866
      11'hdc: T=64'b1101010110011110010011101111111101111000110001111010101110100001;  // -711045377 2026351521
      11'hdd: T=64'b1101010101101110111001000010010001111000101101101111110110100111;  // -714152924 2025258407
      11'hde: T=64'b1101010100111111011111111101101001111000101001100011110100010000;  // -717258790 2024160528
      11'hdf: T=64'b1101010100010000001000100010100001111000100101010110100111011110;  // -720362968 2023057886
      11'he0: T=64'b1101010011100000110010110001010101111000100001001000010000010011;  // -723465451 2021950483
      11'he1: T=64'b1101010010110001011110101010100001111000011100111000101110110010;  // -726566232 2020838322
      11'he2: T=64'b1101010010000010001100001110100101111000011000101000000010111111;  // -729665303 2019721407
      11'he3: T=64'b1101010001010010111011011101111101111000010100010110001100111010;  // -732762657 2018599738
      11'he4: T=64'b1101010000100011101100011001000101111000010000000011001100101000;  // -735858287 2017473320
      11'he5: T=64'b1101001111110100011111000000011101111000001011101111000010001010;  // -738952185 2016342154
      11'he6: T=64'b1101001111000101010011010100011101111000000111011001101101100100;  // -742044345 2015206244
      11'he7: T=64'b1101001110010110001001010101101001111000000011000011001110110111;  // -745134758 2014065591
      11'he8: T=64'b1101001101100111000001000100011001110111111110101011100110001000;  // -748223418 2012920200
      11'he9: T=64'b1101001100110111111010100001001001110111111010010010110011011000;  // -751310318 2011770072
      11'hea: T=64'b1101001100001000110101101100011101110111110101111000110110101001;  // -754395449 2010615209
      11'heb: T=64'b1101001011011001110010100110101101110111110001011101110000000000;  // -757478805 2009455616
      11'hec: T=64'b1101001010101010110001010000010101110111101101000001011111011111;  // -760560379 2008291295
      11'hed: T=64'b1101001001111011110001101001110101110111101000100100000101000111;  // -763640163 2007122247
      11'hee: T=64'b1101001001001100110011110011100101110111100100000101100000111101;  // -766718151 2005948477
      11'hef: T=64'b1101001000011101110111101110001001110111011111100101110011000010;  // -769794334 2004769986
      11'hf0: T=64'b1101000111101110111101011001111001110111011011000100111011011010;  // -772868706 2003586778
      11'hf1: T=64'b1101000111000000000100110111010101110111010110100010111010001000;  // -775941259 2002398856
      11'hf2: T=64'b1101000110010001001110000110111001110111010001111111101111001101;  // -779011986 2001206221
      11'hf3: T=64'b1101000101100010011001001001000001110111001101011011011010101110;  // -782080880 2000008878
      11'hf4: T=64'b1101000100110011100101111110001001110111001000110101111100101100;  // -785147934 1998806828
      11'hf5: T=64'b1101000100000100110100100110110001110111000100001111010101001011;  // -788213140 1997600075
      11'hf6: T=64'b1101000011010110000101000011010001110110111111100111100100001101;  // -791276492 1996388621
      11'hf7: T=64'b1101000010100111010111010100001101110110111010111110101001110110;  // -794337981 1995172470
      11'hf8: T=64'b1101000001111000101011011001111001110110110110010100100110001000;  // -797397602 1993951624
      11'hf9: T=64'b1101000001001010000001010100111001110110110001101001011001000110;  // -800455346 1992726086
      11'hfa: T=64'b1101000000011011011001000101100101110110101100111101000010110011;  // -803511207 1991495859
      11'hfb: T=64'b1100111111101100110010101100100001110110101000001111100011010001;  // -806565176 1990260945
      11'hfc: T=64'b1100111110111110001110001010000001110110100011100000111010100101;  // -809617248 1989021349
      11'hfd: T=64'b1100111110001111101011011110100101110110011110110001001000110000;  // -812667415 1987777072
      11'hfe: T=64'b1100111101100001001010101010101001110110011010000000001101110101;  // -815715670 1986528117
      11'hff: T=64'b1100111100110010101011101110101101110110010101001110001001111000;  // -818762005 1985274488
      11'h100: T=64'b1100111100000100001110101011001101110110010000011010111100111100;  // -821806413 1984016188
      11'h101: T=64'b1100111011010101110011100000100001110110001011100110100111000011;  // -824848888 1982753219
      11'h102: T=64'b1100111010100111011010001111001101110110000110110001001000010000;  // -827889421 1981485584
      11'h103: T=64'b1100111001111001000010110111100101110110000001111010100000100111;  // -830928007 1980213287
      11'h104: T=64'b1100111001001010101101011010001101110101111101000010110000001010;  // -833964637 1978936330
      11'h105: T=64'b1100111000011100011001110111011101110101111000001001110110111100;  // -836999305 1977654716
      11'h106: T=64'b1100110111101110001000001111110101110101110011001111110101000001;  // -840032003 1976368449
      11'h107: T=64'b1100110110111111111000100011101101110101101110010100101010011100;  // -843062725 1975077532
      11'h108: T=64'b1100110110010001101010110011100101110101101001011000010111001110;  // -846091463 1973781966
      11'h109: T=64'b1100110101100011011110111111111001110101100100011010111011011100;  // -849118210 1972481756
      11'h10a: T=64'b1100110100110101010101001001000101110101011111011100010111001001;  // -852142959 1971176905
      11'h10b: T=64'b1100110100000111001101001111100101110101011010011100101010011000;  // -855165703 1969867416
      11'h10c: T=64'b1100110011011001000111010011111001110101010101011011110101001011;  // -858186434 1968553291
      11'h10d: T=64'b1100110010101011000011010110011001110101010000011001110111100110;  // -861205146 1967234534
      11'h10e: T=64'b1100110001111101000001010111100001110101001011010110110001101011;  // -864221832 1965911147
      11'h10f: T=64'b1100110001001111000001010111110001110101000110010010100011011111;  // -867236484 1964583135
      11'h110: T=64'b1100110000100001000011010111100101110101000001001101001101000100;  // -870249095 1963250500
      11'h111: T=64'b1100101111110011000111010111011001110100111100000110101110011110;  // -873259658 1961913246
      11'h112: T=64'b1100101111000101001101010111100101110100110110111111000111101110;  // -876268167 1960571374
      11'h113: T=64'b1100101110010111010101011000101001110100110001110110011000111010;  // -879274614 1959224890
      11'h114: T=64'b1100101101101001011111011011000101110100101100101100100010000011;  // -882278991 1957873795
      11'h115: T=64'b1100101100111011101011011111001101110100100111100001100011001101;  // -885281293 1956518093
      11'h116: T=64'b1100101100001101111001100101100101110100100010010101011100011011;  // -888281511 1955157787
      11'h117: T=64'b1100101011100000001001101110100001110100011101001000001101110000;  // -891279640 1953792880
      11'h118: T=64'b1100101010110010011011111010101001110100010111111001110111010000;  // -894275670 1952423376
      11'h119: T=64'b1100101010000100110000001010001101110100010010101010011000111110;  // -897269597 1951049278
      11'h11a: T=64'b1100101001010111000110011101110001110100001101011001110010111100;  // -900261412 1949670588
      11'h11b: T=64'b1100101000101001011110110101101101110100001000001000000101001111;  // -903251109 1948287311
      11'h11c: T=64'b1100100111111011111001010010011101110100000010110101001111111010;  // -906238681 1946899450
      11'h11d: T=64'b1100100111001110010101110100100001110011111101100001010010111111;  // -909224120 1945507007
      11'h11e: T=64'b1100100110100000110100011100010101110011111000001100001110100010;  // -912207419 1944109986
      11'h11f: T=64'b1100100101110011010101001010010001110011110010110110000010100111;  // -915188572 1942708391
      11'h120: T=64'b1100100101000101110111111110110101110011101101011110101111010000;  // -918167571 1941302224
      11'h121: T=64'b1100100100011000011100111010011001110011101000000110010100100001;  // -921144410 1939891489
      11'h122: T=64'b1100100011101011000011111101011001110011100010101100110010011101;  // -924119082 1938476189
      11'h123: T=64'b1100100010111101101101001000011001110011011101010010001001001000;  // -927091578 1937056328
      11'h124: T=64'b1100100010010000011000011011101001110011010111110110011000100101;  // -930061894 1935631909
      11'h125: T=64'b1100100001100011000101110111110001110011010010011001100000110111;  // -933030020 1934202935
      11'h126: T=64'b1100100000110101110101011101000001110011001100111011100010000010;  // -935995952 1932769410
      11'h127: T=64'b1100100000001000100111001100000001110011000111011100011100001001;  // -938959680 1931331337
      11'h128: T=64'b1100011111011011011011000101000001110011000001111100001111001111;  // -941921200 1929888719
      11'h129: T=64'b1100011110101110010001001000101001110010111100011010111011011000;  // -944880502 1928441560
      11'h12a: T=64'b1100011110000001001001010111001001110010110110111000100000100111;  // -947837582 1926989863
      11'h12b: T=64'b1100011101010100000011110001000101110010110001010100111111000000;  // -950792431 1925533632
      11'h12c: T=64'b1100011100100111000000010110110101110010101011110000010110100110;  // -953745043 1924072870
      11'h12d: T=64'b1100011011111001111111001000111001110010100110001010100111011100;  // -956695410 1922607580
      11'h12e: T=64'b1100011011001101000000000111100101110010100000100011110001100110;  // -959643527 1921137766
      11'h12f: T=64'b1100011010100000000011010011011101110010011010111011110101001000;  // -962589385 1919663432
      11'h130: T=64'b1100011001110011001000101100111001110010010101010010110010000100;  // -965532978 1918184580
      11'h131: T=64'b1100011001000110010000010100010101110010001111101000101000011111;  // -968474299 1916701215
      11'h132: T=64'b1100011000011001011010001010001101110010001001111101011000011011;  // -971413341 1915213339
      11'h133: T=64'b1100010111101100100110001110111001110010000100010001000001111101;  // -974350098 1913720957
      11'h134: T=64'b1100010110111111110100100010111101110001111110100011100101001000;  // -977284561 1912224072
      11'h135: T=64'b1100010110010011000101000110101101110001111000110101000001111111;  // -980216725 1910722687
      11'h136: T=64'b1100010101100110010111111010100101110001110011000101011000100110;  // -983146583 1909216806
      11'h137: T=64'b1100010100111001101100111111000101110001101101010100101001000000;  // -986074127 1907706432
      11'h138: T=64'b1100010100001101000100010100100101110001100111100010110011010001;  // -988999351 1906191569
      11'h139: T=64'b1100010011100000011101111011100101110001100001101111110111011101;  // -991922247 1904672221
      11'h13a: T=64'b1100010010110011111001110100011101110001011011111011110101100111;  // -994842809 1903148391
      11'h13b: T=64'b1100010010000111010111111111100101110001010110000110101101110011;  // -997761031 1901620083
      11'h13c: T=64'b1100010001011010111000011101011101110001010000010000100000000100;  // -1000676905 1900087300
      11'h13d: T=64'b1100010000101110011011001110100101110001001010011001001100011110;  // -1003590423 1898550046
      11'h13e: T=64'b1100010000000010000000010011001101110001000100100000110011000100;  // -1006501581 1897008324
      11'h13f: T=64'b1100001111010101100111101011111001110000111110100111010011111011;  // -1009410370 1895462139
      11'h140: T=64'b1100001110101001010001011001000001110000111000101100101111000101;  // -1012316784 1893911493
      11'h141: T=64'b1100001101111100111101011011000101110000110010110001000100100111;  // -1015220815 1892356391
      11'h142: T=64'b1100001101010000101011110010011001110000101100110100010100100100;  // -1018122458 1890796836
      11'h143: T=64'b1100001100100100011100011111011101110000100110110110011111000000;  // -1021021705 1889232832
      11'h144: T=64'b1100001011111000001111100010101101110000100000110111100011111110;  // -1023918549 1887664382
      11'h145: T=64'b1100001011001100000100111100011101110000011010110111100011100010;  // -1026812985 1886091490
      11'h146: T=64'b1100001010011111111100101101010101110000010100110110011101110000;  // -1029705003 1884514160
      11'h147: T=64'b1100001001110011110110110101100101110000001110110100010010101100;  // -1032594599 1882932396
      11'h148: T=64'b1100001001000111110011010101101101110000001000110001000010011001;  // -1035481765 1881346201
      11'h149: T=64'b1100001000011011110010001110000101110000000010101100101100111011;  // -1038366495 1879755579
      11'h14a: T=64'b1100000111101111110011011111001101101111111100100111010010010110;  // -1041248781 1878160534
      11'h14b: T=64'b1100000111000011110111001001011101101111110110100000110010101101;  // -1044128617 1876561069
      11'h14c: T=64'b1100000110010111111101001101010001101111110000011001001110000100;  // -1047005996 1874957188
      11'h14d: T=64'b1100000101101100000101101011000101101111101010010000100100100000;  // -1049880911 1873348896
      11'h14e: T=64'b1100000101000000010000100011010001101111100100000110110110000011;  // -1052753356 1871736195
      11'h14f: T=64'b1100000100010100011101110110010001101111011101111100000010110010;  // -1055623324 1870119090
      11'h150: T=64'b1100000011101000101101100100100101101111010111110000001010110001;  // -1058490807 1868497585
      11'h151: T=64'b1100000010111100111111101110100001101111010001100011001110000011;  // -1061355800 1866871683
      11'h152: T=64'b1100000010010001010100010100100001101111001011010101001100101011;  // -1064218296 1865241387
      11'h153: T=64'b1100000001100101101011010111000101101111000101000110000110101111;  // -1067078287 1863606703
      11'h154: T=64'b1100000000111010000100110110100101101110111110110101111100010001;  // -1069935767 1861967633
      11'h155: T=64'b1100000000001110100000110011011001101110111000100100101101010110;  // -1072790730 1860324182
      11'h156: T=64'b1011111111100010111111001110000001101110110010010010011010000010;  // -1075643168 1858676354
      11'h157: T=64'b1011111110110111100000000110110101101110101011111111000010011000;  // -1078493075 1857024152
      11'h158: T=64'b1011111110001100000011011110001101101110100101101010100110011100;  // -1081340445 1855367580
      11'h159: T=64'b1011111101100000101001010100101001101110011111010101000110010010;  // -1084185270 1853706642
      11'h15a: T=64'b1011111100110101010001101010100101101110011000111110100001111111;  // -1087027543 1852041343
      11'h15b: T=64'b1011111100001001111100100000010101101110010010100110111001100101;  // -1089867259 1850371685
      11'h15c: T=64'b1011111011011110101001110110011001101110001100001110001101001001;  // -1092704410 1848697673
      11'h15d: T=64'b1011111010110011011001101101001001101110000101110100011100101111;  // -1095538990 1847019311
      11'h15e: T=64'b1011111010001000001100000101000001101101111111011001101000011011;  // -1098370992 1845336603
      11'h15f: T=64'b1011111001011101000000111110011001101101111000111101110000010000;  // -1101200410 1843649552
      11'h160: T=64'b1011111000110001111000011001110001101101110010100000110100010100;  // -1104027236 1841958164
      11'h161: T=64'b1011111000000110110010010111100001101101101100000010110100101000;  // -1106851464 1840262440
      11'h162: T=64'b1011110111011011101110111000000001101101100101100011110001010011;  // -1109673088 1838562387
      11'h163: T=64'b1011110110110000101101111011101101101101011111000011101010010111;  // -1112492101 1836858007
      11'h164: T=64'b1011110110000101101111100011000001101101011000100010011111111001;  // -1115308496 1835149305
      11'h165: T=64'b1011110101011010110011101110011001101101010010000000010001111101;  // -1118122266 1833436285
      11'h166: T=64'b1011110100101111111010011110001001101101001011011101000000100111;  // -1120933406 1831718951
      11'h167: T=64'b1011110100000101000011110010110101101101000100111000101011111010;  // -1123741907 1829997306
      11'h168: T=64'b1011110011011010001111101100101101101100111110010011010011111011;  // -1126547765 1828271355
      11'h169: T=64'b1011110010101111011110001100010001101100110111101100111000101110;  // -1129350972 1826541102
      11'h16a: T=64'b1011110010000100101111010001111101101100110001000101011010010111;  // -1132151521 1824806551
      11'h16b: T=64'b1011110001011010000010111110001001101100101010011100111000111010;  // -1134949406 1823067706
      11'h16c: T=64'b1011110000101111011001010001010001101100100011110011010100011011;  // -1137744620 1821324571
      11'h16d: T=64'b1011110000000100110010001011101101101100011101001000101100111111;  // -1140537157 1819577151
      11'h16e: T=64'b1011101111011010001101101101110101101100010110011101000010101000;  // -1143327011 1817825448
      11'h16f: T=64'b1011101110101111101011111000001001101100001111110000010101011101;  // -1146114174 1816069469
      11'h170: T=64'b1011101110000101001100101011000001101100001001000010100101011111;  // -1148898640 1814309215
      11'h171: T=64'b1011101101011010110000000110110101101100000010010011110010110101;  // -1151680403 1812544693
      11'h172: T=64'b1011101100110000010110001100000101101011111011100011111101100010;  // -1154459455 1810775906
      11'h173: T=64'b1011101100000101111110111011000101101011110100110011000101101001;  // -1157235791 1809002857
      11'h174: T=64'b1011101011011011101010010100010001101011101110000001001011010000;  // -1160009404 1807225552
      11'h175: T=64'b1011101010110001011000011000000001101011100111001110001110011010;  // -1162780288 1805443994
      11'h176: T=64'b1011101010000111001001000110110101101011100000011010001111001100;  // -1165548435 1803658188
      11'h177: T=64'b1011101001011100111100100001000101101011011001100101001101101010;  // -1168313839 1801868138
      11'h178: T=64'b1011101000110010110010100111000101101011010010101111001001111000;  // -1171076495 1800073848
      11'h179: T=64'b1011101000001000101011011001010101101011001011111000000011111010;  // -1173836395 1798275322
      11'h17a: T=64'b1011100111011110100110111000010001101011000100111111111011110100;  // -1176593532 1796472564
      11'h17b: T=64'b1011100110110100100101000100001101101010111110000110110001101011;  // -1179347901 1794665579
      11'h17c: T=64'b1011100110001010100101111101100101101010110111001100100101100100;  // -1182099495 1792854372
      11'h17d: T=64'b1011100101100000101001100100110001101010110000010001010111100001;  // -1184848308 1791038945
      11'h17e: T=64'b1011100100110110101111111010010001101010101001010101000111101000;  // -1187594332 1789219304
      11'h17f: T=64'b1011100100001100111000111110011101101010100010010111110101111101;  // -1190337561 1787395453
      11'h180: T=64'b1011100011100011000100110001101001101010011011011001100010100011;  // -1193077990 1785567395
      11'h181: T=64'b1011100010111001010011010100010101101010010100011010001101100001;  // -1195815611 1783735137
      11'h182: T=64'b1011100010001111100100100110110101101010001101011001110110111000;  // -1198550419 1781898680
      11'h183: T=64'b1011100001100101111000101001101001101010000110011000011110101111;  // -1201282406 1780058031
      11'h184: T=64'b1011100000111100001111011101001001101001111111010110000101001010;  // -1204011566 1778213194
      11'h185: T=64'b1011100000010010101001000001101001101001111000010010101010001100;  // -1206737894 1776364172
      11'h186: T=64'b1011011111101001000101010111101101101001110001001110001101111010;  // -1209461381 1774510970
      11'h187: T=64'b1011011110111111100100011111100101101001101010001000110000011000;  // -1212182023 1772653592
      11'h188: T=64'b1011011110010110000110011001110001101001100011000010010001101011;  // -1214899812 1770792043
      11'h189: T=64'b1011011101101100101011000110100101101001011011111010110001111000;  // -1217614743 1768926328
      11'h18a: T=64'b1011011101000011010010100110100001101001010100110010010001000001;  // -1220326808 1767056449
      11'h18b: T=64'b1011011100011001111100111001111001101001001101101000101111001101;  // -1223036002 1765182413
      11'h18c: T=64'b1011011011110000101010000001001001101001000110011110001100011111;  // -1225742318 1763304223
      11'h18d: T=64'b1011011011000111011001111100101101101000111111010010101000111100;  // -1228445749 1761421884
      11'h18e: T=64'b1011011010011110001100101100111001101000111000000110000100101001;  // -1231146290 1759535401
      11'h18f: T=64'b1011011001110101000010010010001001101000110000111000011111101000;  // -1233843934 1757644776
      11'h190: T=64'b1011011001001011111010101100110101101000101001101001111010000000;  // -1236538675 1755750016
      11'h191: T=64'b1011011000100010110101111101011001101000100010011010010011110101;  // -1239230506 1753851125
      11'h192: T=64'b1011010111111001110100000100001101101000011011001001101101001010;  // -1241919421 1751948106
      11'h193: T=64'b1011010111010000110101000001101101101000010011111000000110000101;  // -1244605413 1750040965
      11'h194: T=64'b1011010110100111111000110110001101101000001100100101011110101010;  // -1247288477 1748129706
      11'h195: T=64'b1011010101111110111111100010001001101000000101010001110110111110;  // -1249968606 1746214334
      11'h196: T=64'b1011010101010110001001000101111101100111111101111101001111000100;  // -1252645793 1744294852
      11'h197: T=64'b1011010100101101010101100001111101100111110110100111100111000010;  // -1255320033 1742371266
      11'h198: T=64'b1011010100000100100100110110100101100111101111010000111110111100;  // -1257991319 1740443580
      11'h199: T=64'b1011010011011011110111000100001101100111100111111001010110110110;  // -1260659645 1738511798
      11'h19a: T=64'b1011010010110011001100001011001101100111100000100000101110110110;  // -1263325005 1736575926
      11'h19b: T=64'b1011010010001010100100001100000101100111011001000111000110111111;  // -1265987391 1734635967
      11'h19c: T=64'b1011010001100001111111000111000101100111010001101100011111010111;  // -1268646799 1732691927
      11'h19d: T=64'b1011010000111001011100111100101001100111001010010000111000000001;  // -1271303222 1730743809
      11'h19e: T=64'b1011010000010000111101101101010001100111000010110100010001000011;  // -1273956652 1728791619
      11'h19f: T=64'b1011001111101000100001011001001001100110111011010110101010100001;  // -1276607086 1726835361
      11'h1a0: T=64'b1011001111000000001000000000110101100110110011111000000100011111;  // -1279254515 1724875039
      11'h1a1: T=64'b1011001110010111110001100100101001100110101100011000011111000011;  // -1281898934 1722910659
      11'h1a2: T=64'b1011001101101111011110000100111101100110100100110111111010010000;  // -1284540337 1720942224
      11'h1a3: T=64'b1011001101000111001101100010001101100110011101010110010110001100;  // -1287178717 1718969740
      11'h1a4: T=64'b1011001100011110111111111100110001100110010101110011110010111011;  // -1289814068 1716993211
      11'h1a5: T=64'b1011001011110110110101010101000001100110001110010000010000100001;  // -1292446384 1715012641
      11'h1a6: T=64'b1011001011001110101101101011011001100110000110101011101111000100;  // -1295075658 1713028036
      11'h1a7: T=64'b1011001010100110101001000000001001100101111111000110001110101000;  // -1297701886 1711039400
      11'h1a8: T=64'b1011001001111110100111010011110101100101110111011111101111010010;  // -1300325059 1709046738
      11'h1a9: T=64'b1011001001010110101000100110101101100101101111111000010001000111;  // -1302945173 1707050055
      11'h1aa: T=64'b1011001000101110101100111001001101100101101000001111110100001010;  // -1305562221 1705049354
      11'h1ab: T=64'b1011001000000110110100001011101101100101100000100110011000100010;  // -1308176197 1703044642
      11'h1ac: T=64'b1011000111011110111110011110100101100101011000111011111110010001;  // -1310787095 1701035921
      11'h1ad: T=64'b1011000110110111001011110010010001100101010001010000100101011111;  // -1313394908 1699023199
      11'h1ae: T=64'b1011000110001111011100000111000101100101001001100100001110001110;  // -1315999631 1697006478
      11'h1af: T=64'b1011000101100111101111011101011101100101000001110110111000100100;  // -1318601257 1694985764
      11'h1b0: T=64'b1011000101000000000101110101110001100100111010001000100100100101;  // -1321199780 1692961061
      11'h1b1: T=64'b1011000100011000011111010000011001100100110010011001010010010111;  // -1323795194 1690932375
      11'h1b2: T=64'b1011000011110000111011101101101101100100101010101001000001111110;  // -1326387493 1688899710
      11'h1b3: T=64'b1011000011001001011011001110000001100100100010110111110011011111;  // -1328976672 1686863071
      11'h1b4: T=64'b1011000010100001111101110001111001100100011011000101100110111111;  // -1331562722 1684822463
      11'h1b5: T=64'b1011000001111010100011011001100001100100010011010010011100100001;  // -1334145640 1682777889
      11'h1b6: T=64'b1011000001010011001100000101011001100100001011011110010100001101;  // -1336725418 1680729357
      11'h1b7: T=64'b1011000000101011110111110101110101100100000011101001001110000101;  // -1339302051 1678676869
      11'h1b8: T=64'b1011000000000100100110101011010001100011111011110011001010001111;  // -1341875532 1676620431
      11'h1b9: T=64'b1010111111011101011000100110000001100011110011111100001000110000;  // -1344445856 1674560048
      11'h1ba: T=64'b1010111110110110001101100110100001100011101100000100001001101100;  // -1347013016 1672495724
      11'h1bb: T=64'b1010111110001111000101101101000101100011100100001011001101001001;  // -1349577007 1670427465
      11'h1bc: T=64'b1010111101101000000000111010001001100011011100010001010011001100;  // -1352137822 1668355276
      11'h1bd: T=64'b1010111101000000111111001110000101100011010100010110011011111000;  // -1354695455 1666279160
      11'h1be: T=64'b1010111100011010000000101001010001100011001100011010100111010100;  // -1357249900 1664199124
      11'h1bf: T=64'b1010111011110011000101001100000001100011000100011101110101100011;  // -1359801152 1662115171
      11'h1c0: T=64'b1010111011001100001100110110110001100010111100100000000110101100;  // -1362349204 1660027308
      11'h1c1: T=64'b1010111010100101010111101001111001100010110100100001011010110010;  // -1364894050 1657935538
      11'h1c2: T=64'b1010111001111110100101100101110001100010101100100001110001111011;  // -1367435684 1655839867
      11'h1c3: T=64'b1010111001010111110110101010101101100010100100100001001100001011;  // -1369974101 1653740299
      11'h1c4: T=64'b1010111000110001001010111001001001100010011100011111101001101000;  // -1372509294 1651636840
      11'h1c5: T=64'b1010111000001010100010010001011101100010010100011101001010010111;  // -1375041257 1649529495
      11'h1c6: T=64'b1010110111100011111100110011111101100010001100011001101110011100;  // -1377569985 1647418268
      11'h1c7: T=64'b1010110110111101011010100001000101100010000100010101010101111101;  // -1380095471 1645303165
      11'h1c8: T=64'b1010110110010110111011011001001001100001111100010000000000111110;  // -1382617710 1643184190
      11'h1c9: T=64'b1010110101110000011111011100100101100001110100001001101111100101;  // -1385136695 1641061349
      11'h1ca: T=64'b1010110101001010000110101011101101100001101100000010100001110110;  // -1387652421 1638934646
      11'h1cb: T=64'b1010110100100011110001000110111001100001100011111010010111110110;  // -1390164882 1636804086
      11'h1cc: T=64'b1010110011111101011110101110100101100001011011110001010001101011;  // -1392674071 1634669675
      11'h1cd: T=64'b1010110011010111001111100011000101100001010011100111001111011001;  // -1395179983 1632531417
      11'h1ce: T=64'b1010110010110001000011100100101101100001001011011100010001000110;  // -1397682613 1630389318
      11'h1cf: T=64'b1010110010001010111010110011111101100001000011010000010110110110;  // -1400181953 1628243382
      11'h1d0: T=64'b1010110001100100110101010001000101100000111011000011100000101111;  // -1402677999 1626093615
      11'h1d1: T=64'b1010110000111110110010111100100001100000110010110101101110110110;  // -1405170744 1623940022
      11'h1d2: T=64'b1010110000011000110011110110100101100000101010100111000001001111;  // -1407660183 1621782607
      11'h1d3: T=64'b1010101111110010110111111111101101100000100010010111011000000000;  // -1410146309 1619621376
      11'h1d4: T=64'b1010101111001100111111011000001101100000011010000110110011001110;  // -1412629117 1617456334
      11'h1d5: T=64'b1010101110100111001010000000011101100000010001110101010010111110;  // -1415108601 1615287486
      11'h1d6: T=64'b1010101110000001010111111000110101100000001001100010110111010101;  // -1417584755 1613114837
      11'h1d7: T=64'b1010101101011011101001000001101101100000000001001111100000011000;  // -1420057573 1610938392
      11'h1d8: T=64'b1010101100110101111101011011011001011111111000111011001110001101;  // -1422527050 1608758157
      11'h1d9: T=64'b1010101100010000010101000110010101011111110000100110000000111000;  // -1424993179 1606574136
      11'h1da: T=64'b1010101011101010110000000010110001011111101000001111111000011110;  // -1427455956 1604386334
      11'h1db: T=64'b1010101011000101001110010001001101011111011111111000110101000101;  // -1429915373 1602194757
      11'h1dc: T=64'b1010101010011111101111110001111001011111010111100000110110110010;  // -1432371426 1599999410
      11'h1dd: T=64'b1010101001111010010100100101010001011111001111000111111101101010;  // -1434824108 1597800298
      11'h1de: T=64'b1010101001010100111100101011101001011111000110101110001001110011;  // -1437273414 1595597427
      11'h1df: T=64'b1010101000101111101000000101011001011110111110010011011011010001;  // -1439719338 1593390801
      11'h1e0: T=64'b1010101000001010010110110010111001011110110101110111110010001001;  // -1442161874 1591180425
      11'h1e1: T=64'b1010100111100101001000110100100001011110101101011011001110100001;  // -1444601016 1588966305
      11'h1e2: T=64'b1010100110111111111110001010100101011110100100111101110000011110;  // -1447036759 1586748446
      11'h1e3: T=64'b1010100110011010110110110101011101011110011100011111011000000110;  // -1449469097 1584526854
      11'h1e4: T=64'b1010100101110101110010110101011101011110010100000000000101011101;  // -1451898025 1582301533
      11'h1e5: T=64'b1010100101010000110010001011000001011110001011011111111000101000;  // -1454323536 1580072488
      11'h1e6: T=64'b1010100100101011110100110110011101011110000010111110110001101110;  // -1456745625 1577839726
      11'h1e7: T=64'b1010100100000110111010111000001001011101111010011100110000110010;  // -1459164286 1575603250
      11'h1e8: T=64'b1010100011100010000100010000011101011101110001111001110101111011;  // -1461579513 1573363067
      11'h1e9: T=64'b1010100010111101010000111111101101011101101001010110000001001110;  // -1463991301 1571119182
      11'h1ea: T=64'b1010100010011000100001000110010001011101100000110001010010110000;  // -1466399644 1568871600
      11'h1eb: T=64'b1010100001110011110100100100011101011101011000001011101010100110;  // -1468804537 1566620326
      11'h1ec: T=64'b1010100001001111001011011010101101011101001111100101001000110110;  // -1471205973 1564365366
      11'h1ed: T=64'b1010100000101010100101101001010001011101000110111101101101100101;  // -1473603948 1562106725
      11'h1ee: T=64'b1010100000000110000011010000100101011100111110010101011000110111;  // -1475998455 1559844407
      11'h1ef: T=64'b1010011111100001100100010000111101011100110101101100001010110100;  // -1478389489 1557578420
      11'h1f0: T=64'b1010011110111101001000101010110001011100101101000010000011011111;  // -1480777044 1555308767
      11'h1f1: T=64'b1010011110011000110000011110011001011100100100010111000010111110;  // -1483161114 1553035454
      11'h1f2: T=64'b1010011101110100011011101100000101011100011011101011001001011000;  // -1485541695 1550758488
      11'h1f3: T=64'b1010011101010000001010010100010001011100010010111110010110101111;  // -1487918780 1548477871
      11'h1f4: T=64'b1010011100101011111100010111010001011100001010010000101011001100;  // -1490292364 1546193612
      11'h1f5: T=64'b1010011100000111110001110101011101011100000001100010000110110010;  // -1492662441 1543905714
      11'h1f6: T=64'b1010011011100011101010101111001101011011111000110010101001100110;  // -1495029005 1541614182
      11'h1f7: T=64'b1010011010111111100111000100110001011011110000000010010011110000;  // -1497392052 1539319024
      11'h1f8: T=64'b1010011010011011100110110110100101011011100111010001000101010011;  // -1499751575 1537020243
      11'h1f9: T=64'b1010011001110111101010000100111101011011011110011110111110010101;  // -1502107569 1534717845
      11'h1fa: T=64'b1010011001010011110000110000001101011011010101101011111110111100;  // -1504460029 1532411836
      11'h1fb: T=64'b1010011000101111111010111000110001011011001100111000000111001110;  // -1506808948 1530102222
      11'h1fc: T=64'b1010011000001100001000011110111001011011000100000011010111001110;  // -1509154322 1527789006
      11'h1fd: T=64'b1010010111101000011001100011000001011010111011001101101111000100;  // -1511496144 1525472196
      11'h1fe: T=64'b1010010111000100101110000101011001011010110010010111001110110100;  // -1513834410 1523151796
      11'h1ff: T=64'b1010010110100001000110000110011101011010101001011111110110100100;  // -1516169113 1520827812
      11'h200: T=64'b1010010101111101100001100110011101011010100000100111100110011001;  // -1518500249 1518500249
      11'h201: T=64'b1010010101011010000000100101110001011010010111101110011110011001;  // -1520827812 1516169113
      11'h202: T=64'b1010010100110110100011000100110001011010001110110100011110101010;  // -1523151796 1513834410
      11'h203: T=64'b1010010100010011001001000011110001011010000101111001100111010000;  // -1525472196 1511496144
      11'h204: T=64'b1010010011101111110010100011001001011001111100111101111000010010;  // -1527789006 1509154322
      11'h205: T=64'b1010010011001100011111100011001001011001110100000001010001110100;  // -1530102222 1506808948
      11'h206: T=64'b1010010010101001010000000100010001011001101011000011110011111101;  // -1532411836 1504460029
      11'h207: T=64'b1010010010000110000100000110101101011001100010000101011110110001;  // -1534717845 1502107569
      11'h208: T=64'b1010010001100010111011101010110101011001011001000110010010010111;  // -1537020243 1499751575
      11'h209: T=64'b1010010000111111110110110001000001011001010000000110001110110100;  // -1539319024 1497392052
      11'h20a: T=64'b1010010000011100110101011001101001011001000111000101010100001101;  // -1541614182 1495029005
      11'h20b: T=64'b1010001111111001110111100100111001011000111110000011100010101001;  // -1543905714 1492662441
      11'h20c: T=64'b1010001111010110111101010011010001011000110101000000111010001100;  // -1546193612 1490292364
      11'h20d: T=64'b1010001110110100000110100101000101011000101011111101011010111100;  // -1548477871 1487918780
      11'h20e: T=64'b1010001110010001010011011010100001011000100010111001000100111111;  // -1550758488 1485541695
      11'h20f: T=64'b1010001101101110100011110100001001011000011001110011111000011010;  // -1553035454 1483161114
      11'h210: T=64'b1010001101001011110111110010000101011000010000101101110101010100;  // -1555308767 1480777044
      11'h211: T=64'b1010001100101001001111010100110001011000000111100110111011110001;  // -1557578420 1478389489
      11'h212: T=64'b1010001100000110101010011100100101010111111110011111001011110111;  // -1559844407 1475998455
      11'h213: T=64'b1010001011100100001001001001101101010111110101010110100101101100;  // -1562106725 1473603948
      11'h214: T=64'b1010001011000001101011011100101001010111101100001101001001010101;  // -1564365366 1471205973
      11'h215: T=64'b1010001010011111010001010101101001010111100011000010110110111001;  // -1566620326 1468804537
      11'h216: T=64'b1010001001111100111010110101000001010111011001110111101110011100;  // -1568871600 1466399644
      11'h217: T=64'b1010001001011010100111111011001001010111010000101011110000000101;  // -1571119182 1463991301
      11'h218: T=64'b1010001000111000011000101000010101010111000111011110111011111001;  // -1573363067 1461579513
      11'h219: T=64'b1010001000010110001100111100111001010110111110010001010001111110;  // -1575603250 1459164286
      11'h21a: T=64'b1010000111110100000100111001001001010110110101000010110010011001;  // -1577839726 1456745625
      11'h21b: T=64'b1010000111010010000000011101100001010110101011110011011101010000;  // -1580072488 1454323536
      11'h21c: T=64'b1010000110101111111111101010001101010110100010100011010010101001;  // -1582301533 1451898025
      11'h21d: T=64'b1010000110001110000010011111101001010110011001010010010010101001;  // -1584526854 1449469097
      11'h21e: T=64'b1010000101101100001000111110001001010110010000000000011101010111;  // -1586748446 1447036759
      11'h21f: T=64'b1010000101001010010011000101111101010110000110101101110010111000;  // -1588966305 1444601016
      11'h220: T=64'b1010000100101000100000110111011101010101111101011010010011010010;  // -1591180425 1442161874
      11'h221: T=64'b1010000100000110110010010010111101010101110100000101111110101010;  // -1593390801 1439719338
      11'h222: T=64'b1010000011100101000111011000110101010101101010110000110101000110;  // -1595597427 1437273414
      11'h223: T=64'b1010000011000011100000001001011001010101100001011010110110101100;  // -1597800298 1434824108
      11'h224: T=64'b1010000010100001111100100100111001010101011000000100000011100010;  // -1599999410 1432371426
      11'h225: T=64'b1010000010000000011100101011101101010101001110101100011011101101;  // -1602194757 1429915373
      11'h226: T=64'b1010000001011111000000011110001001010101000101010011111111010100;  // -1604386334 1427455956
      11'h227: T=64'b1010000000111101100111111100100001010100111011111010101110011011;  // -1606574136 1424993179
      11'h228: T=64'b1010000000011100010011000111001101010100110010100000101001001010;  // -1608758157 1422527050
      11'h229: T=64'b1001111111111011000001111110100001010100101001000101101111100101;  // -1610938392 1420057573
      11'h22a: T=64'b1001111111011001110100100010101101010100011111101010000001110011;  // -1613114837 1417584755
      11'h22b: T=64'b1001111110111000101010110100001001010100010110001101011111111001;  // -1615287486 1415108601
      11'h22c: T=64'b1001111110010111100100110011001001010100001100110000001001111101;  // -1617456334 1412629117
      11'h22d: T=64'b1001111101110110100010100000000001010100000011010010000000000101;  // -1619621376 1410146309
      11'h22e: T=64'b1001111101010101100011111011000101010011111001110011000010010111;  // -1621782607 1407660183
      11'h22f: T=64'b1001111100110100101001000100101001010011110000010011010000111000;  // -1623940022 1405170744
      11'h230: T=64'b1001111100010011110001111101000101010011100110110010101011101111;  // -1626093615 1402677999
      11'h231: T=64'b1001111011110010111110100100101001010011011101010001010011000001;  // -1628243382 1400181953
      11'h232: T=64'b1001111011010010001110111011101001010011010011101111000110110101;  // -1630389318 1397682613
      11'h233: T=64'b1001111010110001100011000010011101010011001010001100000111001111;  // -1632531417 1395179983
      11'h234: T=64'b1001111010010000111010111001010101010011000000101000010100010111;  // -1634669675 1392674071
      11'h235: T=64'b1001111001110000010110100000101001010010110111000011101110010010;  // -1636804086 1390164882
      11'h236: T=64'b1001111001001111110101111000101001010010101101011110010101000101;  // -1638934646 1387652421
      11'h237: T=64'b1001111000101111011001000001101101010010100011111000001000110111;  // -1641061349 1385136695
      11'h238: T=64'b1001111000001110111111111100001001010010011010010001001001101110;  // -1643184190 1382617710
      11'h239: T=64'b1001110111101110101010101000001101010010010000101001010111101111;  // -1645303165 1380095471
      11'h23a: T=64'b1001110111001110011001000110010001010010000111000000110011000001;  // -1647418268 1377569985
      11'h23b: T=64'b1001110110101110001011010110100101010001111101010111011011101001;  // -1649529495 1375041257
      11'h23c: T=64'b1001110110001110000001011001100001010001110011101101010001101110;  // -1651636840 1372509294
      11'h23d: T=64'b1001110101101101111011001111010101010001101010000010010101010101;  // -1653740299 1369974101
      11'h23e: T=64'b1001110101001101111000111000010101010001100000010110100110100100;  // -1655839867 1367435684
      11'h23f: T=64'b1001110100101101111010010100111001010001010110101010000101100010;  // -1657935538 1364894050
      11'h240: T=64'b1001110100001101111111100101010001010001001100111100110010010100;  // -1660027308 1362349204
      11'h241: T=64'b1001110011101110001000101001110101010001000011001110101101000000;  // -1662115171 1359801152
      11'h242: T=64'b1001110011001110010101100010110001010000111001011111110101101100;  // -1664199124 1357249900
      11'h243: T=64'b1001110010101110100110010000100001010000101111110000001100011111;  // -1666279160 1354695455
      11'h244: T=64'b1001110010001110111010110011010001010000100101111111110001011110;  // -1668355276 1352137822
      11'h245: T=64'b1001110001101111010011001011011101010000011100001110100100101111;  // -1670427465 1349577007
      11'h246: T=64'b1001110001001111101111011001010001010000010010011100100110011000;  // -1672495724 1347013016
      11'h247: T=64'b1001110000110000001111011101000001010000001000101001110110100000;  // -1674560048 1344445856
      11'h248: T=64'b1001110000010000110011010111000101001111111110110110010101001100;  // -1676620431 1341875532
      11'h249: T=64'b1001101111110001011011000111101101001111110101000010000010100011;  // -1678676869 1339302051
      11'h24a: T=64'b1001101111010010000110101111001101001111101011001100111110101010;  // -1680729357 1336725418
      11'h24b: T=64'b1001101110110010110110001101111101001111100001010111001001101000;  // -1682777889 1334145640
      11'h24c: T=64'b1001101110010011101001100100000101001111010111100000100011100010;  // -1684822463 1331562722
      11'h24d: T=64'b1001101101110100100000110010000101001111001101101001001100100000;  // -1686863071 1328976672
      11'h24e: T=64'b1001101101010101011011111000001001001111000011110001000100100101;  // -1688899710 1326387493
      11'h24f: T=64'b1001101100110110011010110110100101001110111001111000001011111010;  // -1690932375 1323795194
      11'h250: T=64'b1001101100010111011101101101101101001110101111111110100010100100;  // -1692961061 1321199780
      11'h251: T=64'b1001101011111000100100011101110001001110100110000100001000101001;  // -1694985764 1318601257
      11'h252: T=64'b1001101011011001101111000111001001001110011100001000111110001111;  // -1697006478 1315999631
      11'h253: T=64'b1001101010111010111101101010000101001110010010001101000011011100;  // -1699023199 1313394908
      11'h254: T=64'b1001101010011100010000000110111101001110001000010000011000010111;  // -1701035921 1310787095
      11'h255: T=64'b1001101001111101100110011101111001001101111110010010111101000101;  // -1703044642 1308176197
      11'h256: T=64'b1001101001011111000000101111011001001101110100010100110001101101;  // -1705049354 1305562221
      11'h257: T=64'b1001101001000000011110111011100101001101101010010101110110010101;  // -1707050055 1302945173
      11'h258: T=64'b1001101000100010000001000010111001001101100000010110001011000011;  // -1709046738 1300325059
      11'h259: T=64'b1001101000000011100111000101100001001101010110010101101111111110;  // -1711039400 1297701886
      11'h25a: T=64'b1001100111100101010001000011110001001101001100010100100101001010;  // -1713028036 1295075658
      11'h25b: T=64'b1001100111000110111110111101111101001101000010010010101010110000;  // -1715012641 1292446384
      11'h25c: T=64'b1001100110101000110000110100010101001100111000010000000000110100;  // -1716993211 1289814068
      11'h25d: T=64'b1001100110001010100110100111010001001100101110001100100111011101;  // -1718969740 1287178717
      11'h25e: T=64'b1001100101101100100000010111000001001100100100001000011110110001;  // -1720942224 1284540337
      11'h25f: T=64'b1001100101001110011110000011110101001100011010000011100110110110;  // -1722910659 1281898934
      11'h260: T=64'b1001100100110000011111101110000101001100001111111101111111110011;  // -1724875039 1279254515
      11'h261: T=64'b1001100100010010100101010101111101001100000101110111101001101110;  // -1726835361 1276607086
      11'h262: T=64'b1001100011110100101110111011110101001011111011110000100100101100;  // -1728791619 1273956652
      11'h263: T=64'b1001100011010110111100011111111101001011110001101000110000110110;  // -1730743809 1271303222
      11'h264: T=64'b1001100010111001001110000010100101001011100111100000001110001111;  // -1732691927 1268646799
      11'h265: T=64'b1001100010011011100011100100000101001011011101010110111100111111;  // -1734635967 1265987391
      11'h266: T=64'b1001100001111101111101000100101001001011010011001100111101001101;  // -1736575926 1263325005
      11'h267: T=64'b1001100001100000011010100100101001001011001001000010001110111101;  // -1738511798 1260659645
      11'h268: T=64'b1001100001000010111100000100010001001010111110110110110010010111;  // -1740443580 1257991319
      11'h269: T=64'b1001100000100101100001100011111001001010110100101010100111100001;  // -1742371266 1255320033
      11'h26a: T=64'b1001100000001000001011000011110001001010101010011101101110100001;  // -1744294852 1252645793
      11'h26b: T=64'b1001011111101010111000100100001001001010100000010000000111011110;  // -1746214334 1249968606
      11'h26c: T=64'b1001011111001101101010000101011001001010010110000001110010011101;  // -1748129706 1247288477
      11'h26d: T=64'b1001011110110000011111100111101101001010001011110010101111100101;  // -1750040965 1244605413
      11'h26e: T=64'b1001011110010011011001001011011001001010000001100010111110111101;  // -1751948106 1241919421
      11'h26f: T=64'b1001011101110110010110110000101101001001110111010010100000101010;  // -1753851125 1239230506
      11'h270: T=64'b1001011101011001011000011000000001001001101101000001010100110011;  // -1755750016 1236538675
      11'h271: T=64'b1001011100111100011110000001100001001001100010101111011011011110;  // -1757644776 1233843934
      11'h272: T=64'b1001011100011111100111101101011101001001011000011100110100110010;  // -1759535401 1231146290
      11'h273: T=64'b1001011100000010110101011100010001001001001110001001100000110101;  // -1761421884 1228445749
      11'h274: T=64'b1001011011100110000111001110000101001001000011110101011111101110;  // -1763304223 1225742318
      11'h275: T=64'b1001011011001001011101000011001101001000111001100000110001100010;  // -1765182413 1223036002
      11'h276: T=64'b1001011010101100110110111011111101001000101111001011010110011000;  // -1767056449 1220326808
      11'h277: T=64'b1001011010010000010100111000100001001000100100110101001110010111;  // -1768926328 1217614743
      11'h278: T=64'b1001011001110011110110111001010101001000011010011110011001100100;  // -1770792043 1214899812
      11'h279: T=64'b1001011001010111011100111110100001001000010000000110111000000111;  // -1772653592 1212182023
      11'h27a: T=64'b1001011000111011000111001000011001001000000101101110101010000101;  // -1774510970 1209461381
      11'h27b: T=64'b1001011000011110110101010111010001000111111011010101101111100110;  // -1776364172 1206737894
      11'h27c: T=64'b1001011000000010100111101011011001000111110000111100001000101110;  // -1778213194 1204011566
      11'h27d: T=64'b1001010111100110011110000101000101000111100110100001110101100110;  // -1780058031 1201282406
      11'h27e: T=64'b1001010111001010011000100100100001000111011100000110110110010011;  // -1781898680 1198550419
      11'h27f: T=64'b1001010110101110010111001001111101000111010001101011001010111011;  // -1783735137 1195815611
      11'h280: T=64'b1001010110010010011001110101110101000111000111001110110011100110;  // -1785567395 1193077990
      11'h281: T=64'b1001010101110110100000101000001101000110111100110001110000011001;  // -1787395453 1190337561
      11'h282: T=64'b1001010101011010101011100001100001000110110010010100000001011100;  // -1789219304 1187594332
      11'h283: T=64'b1001010100111110111010100001111101000110100111110101100110110100;  // -1791038945 1184848308
      11'h284: T=64'b1001010100100011001101101001110001000110011101010110100000100111;  // -1792854372 1182099495
      11'h285: T=64'b1001010100000111100100111001010101000110010010110110101110111101;  // -1794665579 1179347901
      11'h286: T=64'b1001010011101100000000010000110001000110001000010110010001111100;  // -1796472564 1176593532
      11'h287: T=64'b1001010011010000011111110000011001000101111101110101001001101011;  // -1798275322 1173836395
      11'h288: T=64'b1001010010110101000011011000100001000101110011010011010110001111;  // -1800073848 1171076495
      11'h289: T=64'b1001010010011001101011001001011001000101101000110000110111101111;  // -1801868138 1168313839
      11'h28a: T=64'b1001010001111110010111000011010001000101011110001101101110010011;  // -1803658188 1165548435
      11'h28b: T=64'b1001010001100011000111000110011001000101010011101001111010000000;  // -1805443994 1162780288
      11'h28c: T=64'b1001010001000111111011010011000001000101001001000101011010111100;  // -1807225552 1160009404
      11'h28d: T=64'b1001010000101100110011101001011101000100111110100000010001001111;  // -1809002857 1157235791
      11'h28e: T=64'b1001010000010001110000001001111001000100110011111010011100111111;  // -1810775906 1154459455
      11'h28f: T=64'b1001001111110110110000110100101101000100101001010011111110010011;  // -1812544693 1151680403
      11'h290: T=64'b1001001111011011110101101010000101000100011110101100110101010000;  // -1814309215 1148898640
      11'h291: T=64'b1001001111000000111110101010001101000100010100000101000001111110;  // -1816069469 1146114174
      11'h292: T=64'b1001001110100110001011110101100001000100001001011100100100100011;  // -1817825448 1143327011
      11'h293: T=64'b1001001110001011011101001100000101000011111110110011011101000101;  // -1819577151 1140537157
      11'h294: T=64'b1001001101110000110010101110010101000011110100001001101011101100;  // -1821324571 1137744620
      11'h295: T=64'b1001001101010110001100011100011001000011101001011111010000011110;  // -1823067706 1134949406
      11'h296: T=64'b1001001100111011101010010110100101000011011110110100001011100001;  // -1824806551 1132151521
      11'h297: T=64'b1001001100100001001100011101001001000011010100001000011100111100;  // -1826541102 1129350972
      11'h298: T=64'b1001001100000110110010110000010101000011001001011100000100110101;  // -1828271355 1126547765
      11'h299: T=64'b1001001011101100011101010000011001000010111110101111000011010011;  // -1829997306 1123741907
      11'h29a: T=64'b1001001011010010001011111101100101000010110100000001011000011110;  // -1831718951 1120933406
      11'h29b: T=64'b1001001010110111111110111000001101000010101001010011000100011010;  // -1833436285 1118122266
      11'h29c: T=64'b1001001010011101110110000000011101000010011110100100000111010000;  // -1835149305 1115308496
      11'h29d: T=64'b1001001010000011110001010110100101000010010011110100100001000101;  // -1836858007 1112492101
      11'h29e: T=64'b1001001001101001110000111010110101000010001001000100010010000000;  // -1838562387 1109673088
      11'h29f: T=64'b1001001001001111110100101101100001000001111110010011011010001000;  // -1840262440 1106851464
      11'h2a0: T=64'b1001001000110101111100101110110001000001110011100001111001100100;  // -1841958164 1104027236
      11'h2a1: T=64'b1001001000011100001000111111000001000001101000101111110000011010;  // -1843649552 1101200410
      11'h2a2: T=64'b1001001000000010011001011110010101000001011101111100111110110000;  // -1845336603 1098370992
      11'h2a3: T=64'b1001000111101000101110001101000101000001010011001001100100101110;  // -1847019311 1095538990
      11'h2a4: T=64'b1001000111001111000111001011011101000001001000010101100010011010;  // -1848697673 1092704410
      11'h2a5: T=64'b1001000110110101100100011001101101000000111101100000110111111011;  // -1850371685 1089867259
      11'h2a6: T=64'b1001000110011100000101111000000101000000110010101011100101010111;  // -1852041343 1087027543
      11'h2a7: T=64'b1001000110000010101011100110111001000000100111110101101010110110;  // -1853706642 1084185270
      11'h2a8: T=64'b1001000101101001010101100110010001000000011100111111001000011101;  // -1855367580 1081340445
      11'h2a9: T=64'b1001000101010000000011110110100001000000010010000111111110010011;  // -1857024152 1078493075
      11'h2aa: T=64'b1001000100110110110110010111111001000000000111010000001100100000;  // -1858676354 1075643168
      11'h2ab: T=64'b1001000100011101101101001010101000111111111100010111110011001010;  // -1860324182 1072790730
      11'h2ac: T=64'b1001000100000100101000001110111100111111110001011110110010010111;  // -1861967633 1069935767
      11'h2ad: T=64'b1001000011101011100111100101000100111111100110100101001010001111;  // -1863606703 1067078287
      11'h2ae: T=64'b1001000011010010101011001101010100111111011011101010111010111000;  // -1865241387 1064218296
      11'h2af: T=64'b1001000010111001110011000111110100111111010000110000000100011000;  // -1866871683 1061355800
      11'h2b0: T=64'b1001000010100000111111010100111100111111000101110100100110110111;  // -1868497585 1058490807
      11'h2b1: T=64'b1001000010001000001111110100111000111110111010111000100010011100;  // -1870119090 1055623324
      11'h2b2: T=64'b1001000001101111100100100111110100111110101111111011110111001100;  // -1871736195 1052753356
      11'h2b3: T=64'b1001000001010110111101101110000000111110100100111110100101001111;  // -1873348896 1049880911
      11'h2b4: T=64'b1001000000111110011011000111110000111110011010000000101100101100;  // -1874957188 1047005996
      11'h2b5: T=64'b1001000000100101111100110101001100111110001111000010001101101001;  // -1876561069 1044128617
      11'h2b6: T=64'b1001000000001101100010110110101000111110000100000011001000001101;  // -1878160534 1041248781
      11'h2b7: T=64'b1000111111110101001101001100010100111101111001000011011100011111;  // -1879755579 1038366495
      11'h2b8: T=64'b1000111111011100111011110110011100111101101110000011001010100101;  // -1881346201 1035481765
      11'h2b9: T=64'b1000111111000100101110110101010000111101100011000010010010100111;  // -1882932396 1032594599
      11'h2ba: T=64'b1000111110101100100110001001000000111101011000000000110100101011;  // -1884514160 1029705003
      11'h2bb: T=64'b1000111110010100100001110001111000111101001100111110110000111001;  // -1886091490 1026812985
      11'h2bc: T=64'b1000111101111100100001110000001000111101000001111100000111010101;  // -1887664382 1023918549
      11'h2bd: T=64'b1000111101100100100110000100000000111100110110111000111000001001;  // -1889232832 1021021705
      11'h2be: T=64'b1000111101001100101110101101110000111100101011110101000011011010;  // -1890796836 1018122458
      11'h2bf: T=64'b1000111100110100111011101101100100111100100000110000101001001111;  // -1892356391 1015220815
      11'h2c0: T=64'b1000111100011101001101000011101100111100010101101011101001110000;  // -1893911493 1012316784
      11'h2c1: T=64'b1000111100000101100010110000010100111100001010100110000101000010;  // -1895462139 1009410370
      11'h2c2: T=64'b1000111011101101111100110011110000111011111111011111111011001101;  // -1897008324 1006501581
      11'h2c3: T=64'b1000111011010110011011001110001000111011110100011001001100010111;  // -1898550046 1003590423
      11'h2c4: T=64'b1000111010111110111101111111110000111011101001010001111000101001;  // -1900087300 1000676905
      11'h2c5: T=64'b1000111010100111100101001000110100111011011110001010000000000111;  // -1901620083 997761031
      11'h2c6: T=64'b1000111010010000010000101001100100111011010011000001100010111001;  // -1903148391 994842809
      11'h2c7: T=64'b1000111001111001000000100010001100111011000111111000100001000111;  // -1904672221 991922247
      11'h2c8: T=64'b1000111001100001110100110010111100111010111100101110111010110111;  // -1906191569 988999351
      11'h2c9: T=64'b1000111001001010101101011100000000111010110001100100110000001111;  // -1907706432 986074127
      11'h2ca: T=64'b1000111000110011101010011101101000111010100110011010000001010111;  // -1909216806 983146583
      11'h2cb: T=64'b1000111000011100101011111000000100111010011011001110101110010101;  // -1910722687 980216725
      11'h2cc: T=64'b1000111000000101110001101011100000111010010000000010110111010001;  // -1912224072 977284561
      11'h2cd: T=64'b1000110111101110111011111000001100111010000100110110011100010010;  // -1913720957 974350098
      11'h2ce: T=64'b1000110111011000001010011110010100111001111001101001011101011101;  // -1915213339 971413341
      11'h2cf: T=64'b1000110111000001011101011110000100111001101110011011111010111011;  // -1916701215 968474299
      11'h2d0: T=64'b1000110110101010110100110111110000111001100011001101110100110010;  // -1918184580 965532978
      11'h2d1: T=64'b1000110110010100010000101011100000111001010111111111001011001001;  // -1919663432 962589385
      11'h2d2: T=64'b1000110101111101110000111001101000111001001100101111111110000111;  // -1921137766 959643527
      11'h2d3: T=64'b1000110101100111010101100010010000111001000001100000001101110010;  // -1922607580 956695410
      11'h2d4: T=64'b1000110101010000111110100101101000111000110110001111111010010011;  // -1924072870 953745043
      11'h2d5: T=64'b1000110100111010101100000100000000111000101010111111000011101111;  // -1925533632 950792431
      11'h2d6: T=64'b1000110100100100011101111101100100111000011111101101101010001110;  // -1926989863 947837582
      11'h2d7: T=64'b1000110100001110010100010010100000111000010100011011101101110110;  // -1928441560 944880502
      11'h2d8: T=64'b1000110011111000001111000011000100111000001001001001001110110000;  // -1929888719 941921200
      11'h2d9: T=64'b1000110011100010001110001111011100110111111101110110001101000000;  // -1931331337 938959680
      11'h2da: T=64'b1000110011001100010001110111111000110111110010100010101000110000;  // -1932769410 935995952
      11'h2db: T=64'b1000110010110110011001111100100100110111100111001110100010000100;  // -1934202935 933030020
      11'h2dc: T=64'b1000110010100000100110011101101100110111011011111001111001000110;  // -1935631909 930061894
      11'h2dd: T=64'b1000110010001010110111011011100000110111010000100100101101111010;  // -1937056328 927091578
      11'h2de: T=64'b1000110001110101001100110110001100110111000101001111000000101010;  // -1938476189 924119082
      11'h2df: T=64'b1000110001011111100110101101111100110110111001111000110001011010;  // -1939891489 921144410
      11'h2e0: T=64'b1000110001001010000101000011000000110110101110100010000000010011;  // -1941302224 918167571
      11'h2e1: T=64'b1000110000110100100111110101100100110110100011001010101101011100;  // -1942708391 915188572
      11'h2e2: T=64'b1000110000011111001111000101111000110110010111110010111000111011;  // -1944109986 912207419
      11'h2e3: T=64'b1000110000001001111010110100000100110110001100011010100010111000;  // -1945507007 909224120
      11'h2e4: T=64'b1000101111110100101011000000011000110110000001000001101011011001;  // -1946899450 906238681
      11'h2e5: T=64'b1000101111011111011111101011000100110101110101101000010010100101;  // -1948287311 903251109
      11'h2e6: T=64'b1000101111001010011000110100010000110101101010001110011000100100;  // -1949670588 900261412
      11'h2e7: T=64'b1000101110110101010110011100001000110101011110110011111101011101;  // -1951049278 897269597
      11'h2e8: T=64'b1000101110100000011000100011000000110101010011011001000001010110;  // -1952423376 894275670
      11'h2e9: T=64'b1000101110001011011111001001000000110101000111111101100100011000;  // -1953792880 891279640
      11'h2ea: T=64'b1000101101110110101010001110010100110100111100100001100110100111;  // -1955157787 888281511
      11'h2eb: T=64'b1000101101100001111001110011001100110100110001000101001000001101;  // -1956518093 885281293
      11'h2ec: T=64'b1000101101001101001101110111110100110100100101101000001001001111;  // -1957873795 882278991
      11'h2ed: T=64'b1000101100111000100110011100011000110100011010001010101001110110;  // -1959224890 879274614
      11'h2ee: T=64'b1000101100100100000011100001001000110100001110101100101010000111;  // -1960571374 876268167
      11'h2ef: T=64'b1000101100001111100101000110001000110100000011001110001010001010;  // -1961913246 873259658
      11'h2f0: T=64'b1000101011111011001011001011110000110011110111101111001010000111;  // -1963250500 870249095
      11'h2f1: T=64'b1000101011100110110101110010000100110011101100001111101010000100;  // -1964583135 867236484
      11'h2f2: T=64'b1000101011010010100100111001010100110011100000101111101010001000;  // -1965911147 864221832
      11'h2f3: T=64'b1000101010111110011000100001101000110011010101001111001010011010;  // -1967234534 861205146
      11'h2f4: T=64'b1000101010101010010000101011010100110011001001101110001011000010;  // -1968553291 858186434
      11'h2f5: T=64'b1000101010010110001101010110100000110010111110001100101100000111;  // -1969867416 855165703
      11'h2f6: T=64'b1000101010000010001110100011011100110010110010101010101101101111;  // -1971176905 852142959
      11'h2f7: T=64'b1000101001101110010100010010010000110010100111001000010000000010;  // -1972481756 849118210
      11'h2f8: T=64'b1000101001011010011110100011001000110010011011100101010011000111;  // -1973781966 846091463
      11'h2f9: T=64'b1000101001000110101101010110010000110010010000000001110111000101;  // -1975077532 843062725
      11'h2fa: T=64'b1000101000110011000000101011111100110010000100011101111100000011;  // -1976368449 840032003
      11'h2fb: T=64'b1000101000011111011000100100010000110001111000111001100010001001;  // -1977654716 836999305
      11'h2fc: T=64'b1000101000001011110100111111011000110001101101010100101001011101;  // -1978936330 833964637
      11'h2fd: T=64'b1000100111111000010101111101100100110001100001101111010010000111;  // -1980213287 830928007
      11'h2fe: T=64'b1000100111100100111011011111000000110001010110001001011100001101;  // -1981485584 827889421
      11'h2ff: T=64'b1000100111010001100101100011110100110001001010100011000111111000;  // -1982753219 824848888
      11'h300: T=64'b1000100110111110010100001100010000110000111110111100010101001101;  // -1984016188 821806413
      11'h301: T=64'b1000100110101011000111011000100000110000110011010101000100010101;  // -1985274488 818762005
      11'h302: T=64'b1000100110010111111111001000101100110000100111101101010101010110;  // -1986528117 815715670
      11'h303: T=64'b1000100110000100111011011101000000110000011100000101001000010111;  // -1987777072 812667415
      11'h304: T=64'b1000100101110001111100010101101100110000010000011100011101100000;  // -1989021349 809617248
      11'h305: T=64'b1000100101011111000001110010111100110000000100110011010100111000;  // -1990260945 806565176
      11'h306: T=64'b1000100101001100001011110100110100101111111001001001101110100111;  // -1991495859 803511207
      11'h307: T=64'b1000100100111001011010011011101000101111101101011111101010110010;  // -1992726086 800455346
      11'h308: T=64'b1000100100100110101101100111100000101111100001110101001001100010;  // -1993951624 797397602
      11'h309: T=64'b1000100100010100000101011000101000101111010110001010001010111101;  // -1995172470 794337981
      11'h30a: T=64'b1000100100000001100001101111001100101111001010011110101111001100;  // -1996388621 791276492
      11'h30b: T=64'b1000100011101111000010101011010100101110111110110010110110010100;  // -1997600075 788213140
      11'h30c: T=64'b1000100011011100101000001101010000101110110011000110100000011110;  // -1998806828 785147934
      11'h30d: T=64'b1000100011001010010010010101001000101110100111011001101101110000;  // -2000008878 782080880
      11'h30e: T=64'b1000100010111000000001000011001100101110011011101100011110010010;  // -2001206221 779011986
      11'h30f: T=64'b1000100010100101110100010111100000101110001111111110110010001011;  // -2002398856 775941259
      11'h310: T=64'b1000100010010011101100010010011000101110000100010000101001100010;  // -2003586778 772868706
      11'h311: T=64'b1000100010000001101000110011111000101101111000100010000100011110;  // -2004769986 769794334
      11'h312: T=64'b1000100001101111101001111100001100101101101100110011000011000111;  // -2005948477 766718151
      11'h313: T=64'b1000100001011101101111101011100100101101100001000011100101100011;  // -2007122247 763640163
      11'h314: T=64'b1000100001001011111010000010000100101101010101010011101011111011;  // -2008291295 760560379
      11'h315: T=64'b1000100000111010001001000000000000101101001001100011010110010101;  // -2009455616 757478805
      11'h316: T=64'b1000100000101000011100100101011100101100111101110010100100111001;  // -2010615209 754395449
      11'h317: T=64'b1000100000010110110100110010100000101100110010000001010111101110;  // -2011770072 751310318
      11'h318: T=64'b1000100000000101010001100111100000101100100110001111101110111010;  // -2012920200 748223418
      11'h319: T=64'b1000011111110011110011000100100100101100011010011101101010100110;  // -2014065591 745134758
      11'h31a: T=64'b1000011111100010011001001001110000101100001110101011001010111001;  // -2015206244 742044345
      11'h31b: T=64'b1000011111010001000011110111011000101100000010111000001111111001;  // -2016342154 738952185
      11'h31c: T=64'b1000011110111111110011001101100000101011110111000100111001101111;  // -2017473320 735858287
      11'h31d: T=64'b1000011110101110100111001100011000101011101011010001001000100001;  // -2018599738 732762657
      11'h31e: T=64'b1000011110011101011111110100000100101011011111011100111100010111;  // -2019721407 729665303
      11'h31f: T=64'b1000011110001100011101000100111000101011010011101000010101011000;  // -2020838322 726566232
      11'h320: T=64'b1000011101111011011110111110110100101011000111110011010011101011;  // -2021950483 723465451
      11'h321: T=64'b1000011101101010100101100010001000101010111011111101110111011000;  // -2023057886 720362968
      11'h322: T=64'b1000011101011001110000101111000000101010110000001000000000100110;  // -2024160528 717258790
      11'h323: T=64'b1000011101001001000000100101100100101010100100010001101111011100;  // -2025258407 714152924
      11'h324: T=64'b1000011100111000010101000101111100101010011000011011000100000001;  // -2026351521 711045377
      11'h325: T=64'b1000011100100111101110010000011000101010001100100011111110011101;  // -2027439866 707936157
      11'h326: T=64'b1000011100010111001100000100111100101010000000101100011110111000;  // -2028523441 704825272
      11'h327: T=64'b1000011100000110101110100011111000101001110100110100100101011000;  // -2029602242 701712728
      11'h328: T=64'b1000011011110110010101101101010000101001101000111100010010000101;  // -2030676268 698598533
      11'h329: T=64'b1000011011100110000001100001010100101001011101000011100101000110;  // -2031745515 695482694
      11'h32a: T=64'b1000011011010101110010000000001100101001010001001010011110100010;  // -2032809981 692365218
      11'h32b: T=64'b1000011011000101100111001010000000101001000101010000111110100001;  // -2033869664 689246113
      11'h32c: T=64'b1000011010110101100000111110111100101000111001010111000101001010;  // -2034924561 686125386
      11'h32d: T=64'b1000011010100101011111011111001100101000101101011100110010100101;  // -2035974669 683003045
      11'h32e: T=64'b1000011010010101100010101010110100101000100001100010000110111001;  // -2037019987 679879097
      11'h32f: T=64'b1000011010000101101010100010000000101000010101100111000010001101;  // -2038060512 676753549
      11'h330: T=64'b1000011001110101110111000101000000101000001001101011100100101000;  // -2039096240 673626408
      11'h331: T=64'b1000011001100110001000010011110100100111111101101111101110010010;  // -2040127171 670497682
      11'h332: T=64'b1000011001010110011110001110101100100111110001110011011111010011;  // -2041153301 667367379
      11'h333: T=64'b1000011001000110111000110101110100100111100101110110110111110001;  // -2042174627 664235505
      11'h334: T=64'b1000011000110111011000001001001100100111011001111001110111110100;  // -2043191149 661102068
      11'h335: T=64'b1000011000100111111100001001001000100111001101111100011111100011;  // -2044202862 657967075
      11'h336: T=64'b1000011000011000100100110101101000100111000001111110101111000110;  // -2045209766 654830534
      11'h337: T=64'b1000011000001001010010001111000000100110110110000000100110100101;  // -2046211856 651692453
      11'h338: T=64'b1000010111111010000100010101010000100110101010000010000110000101;  // -2047209132 648552837
      11'h339: T=64'b1000010111101010111011001000100100100110011110000011001101110000;  // -2048201591 645411696
      11'h33a: T=64'b1000010111011011110110101001001000100110010010000011111101101100;  // -2049189230 642269036
      11'h33b: T=64'b1000010111001100110110110111000100100110000110000100010110000001;  // -2050172047 639124865
      11'h33c: T=64'b1000010110111101111011110010100000100101111010000100010110110110;  // -2051150040 635979190
      11'h33d: T=64'b1000010110101111000101011011101000100101101110000100000000010010;  // -2052123206 632832018
      11'h33e: T=64'b1000010110100000010011110010100100100101100010000011010010011101;  // -2053091543 629683357
      11'h33f: T=64'b1000010110010001100110110111011100100101010110000010001101011110;  // -2054055049 626533214
      11'h340: T=64'b1000010110000010111110101010011000100101001010000000110001011101;  // -2055013722 623381597
      11'h341: T=64'b1000010101110100011011001011100100100100111101111110111110100010;  // -2055967559 620228514
      11'h342: T=64'b1000010101100101111100011011000100100100110001111100110100110010;  // -2056916559 617073970
      11'h343: T=64'b1000010101010111100010011001001000100100100101111010010100010111;  // -2057860718 613917975
      11'h344: T=64'b1000010101001001001101000101110100100100011001110111011101010111;  // -2058800035 610760535
      11'h345: T=64'b1000010100111010111100100001010100100100001101110100001111111010;  // -2059734507 607601658
      11'h346: T=64'b1000010100101100110000101011110000100100000001110000101100000111;  // -2060664132 604441351
      11'h347: T=64'b1000010100011110101001100101001100100011110101101100110010000110;  // -2061588909 601279622
      11'h348: T=64'b1000010100010000100111001101110100100011101001101000100001111110;  // -2062508835 598116478
      11'h349: T=64'b1000010100000010101001100101110100100011011101100011111011110111;  // -2063423907 594951927
      11'h34a: T=64'b1000010011110100110000101101010100100011010001011110111111111000;  // -2064334123 591785976
      11'h34b: T=64'b1000010011100110111100100100010100100011000101011001101110001000;  // -2065239483 588618632
      11'h34c: T=64'b1000010011011001001101001011001000100010111001010100000110101111;  // -2066139982 585449903
      11'h34d: T=64'b1000010011001011100010100001110000100010101101001110001001110100;  // -2067035620 582279796
      11'h34e: T=64'b1000010010111101111100101000011100100010100001000111110111011111;  // -2067926393 579108319
      11'h34f: T=64'b1000010010110000011011011111001100100010010101000001001111111000;  // -2068812301 575935480
      11'h350: T=64'b1000010010100010111111000110001100100010001000111010010011000101;  // -2069693341 572761285
      11'h351: T=64'b1000010010010101100111011101101000100001111100110011000001001111;  // -2070569510 569585743
      11'h352: T=64'b1000010010001000010100100101100100100001110000101011011010011100;  // -2071440807 566408860
      11'h353: T=64'b1000010001111011000110011110001000100001100100100011011110110100;  // -2072307230 563230644
      11'h354: T=64'b1000010001101101111101000111100000100001011000011011001110011111;  // -2073168776 560051103
      11'h355: T=64'b1000010001100000111000100001101100100001001100010010101001100101;  // -2074025445 556870245
      11'h356: T=64'b1000010001010011111000101101000000100001000000001001110000001100;  // -2074877232 553688076
      11'h357: T=64'b1000010001000110111101101001011000100000110100000000100010011100;  // -2075724138 550504604
      11'h358: T=64'b1000010000111010000111010111000100100000100111110111000000011100;  // -2076566159 547319836
      11'h359: T=64'b1000010000101101010101110110001100100000011011101101001010010101;  // -2077403293 544133781
      11'h35a: T=64'b1000010000100000101001000110110100100000001111100011000000001101;  // -2078235539 540946445
      11'h35b: T=64'b1000010000010100000001001001000100100000000011011000100010001101;  // -2079062895 537757837
      11'h35c: T=64'b1000010000000111011101111101000100011111110111001101110000011011;  // -2079885359 534567963
      11'h35d: T=64'b1000001111111010111111100010111100011111101011000010101010111111;  // -2080702929 531376831
      11'h35e: T=64'b1000001111101110100101111010111000011111011110110111010010000000;  // -2081515602 528184448
      11'h35f: T=64'b1000001111100010010001000100111000011111010010101011100101100111;  // -2082323378 524990823
      11'h360: T=64'b1000001111010110000001000001001100011111000110011111100101111011;  // -2083126253 521795963
      11'h361: T=64'b1000001111001001110101101111110100011110111010010011010011000011;  // -2083924227 518599875
      11'h362: T=64'b1000001110111101101111010000111100011110101110000110101101000110;  // -2084717297 515402566
      11'h363: T=64'b1000001110110001101101100100101000011110100001111001110100001101;  // -2085505462 512204045
      11'h364: T=64'b1000001110100101110000101011000100011110010101101100101000011110;  // -2086288719 509004318
      11'h365: T=64'b1000001110011001111000100100010100011110001001011111001010000001;  // -2087067067 505803393
      11'h366: T=64'b1000001110001110000101010000100000011101111101010001011000111111;  // -2087840504 502601279
      11'h367: T=64'b1000001110000010010110101111110000011101110001000011010101011101;  // -2088609028 499397981
      11'h368: T=64'b1000001101110110101101000010001100011101100100110100111111100101;  // -2089372637 496193509
      11'h369: T=64'b1000001101101011001000000111111000011101011000100110010111011101;  // -2090131330 492987869
      11'h36a: T=64'b1000001101011111101000000001000000011101001100010111011101001101;  // -2090885104 489781069
      11'h36b: T=64'b1000001101010100001100101101100100011101000000001000010000111100;  // -2091633959 486573116
      11'h36c: T=64'b1000001101001000110110001101110100011100110011111000110010110011;  // -2092377891 483364019
      11'h36d: T=64'b1000001100111101100100100001110000011100100111101001000010111000;  // -2093116900 480153784
      11'h36e: T=64'b1000001100110010010111101001100000011100011011011001000001010011;  // -2093850984 476942419
      11'h36f: T=64'b1000001100100111001111100101001100011100001111001000101110001100;  // -2094580141 473729932
      11'h370: T=64'b1000001100011100001100010100111100011100000010111000001001101010;  // -2095304369 470516330
      11'h371: T=64'b1000001100010001001101111000111000011011110110100111010011110101;  // -2096023666 467301621
      11'h372: T=64'b1000001100000110010100010001000100011011101010010110001100110101;  // -2096738031 464085813
      11'h373: T=64'b1000001011111011011111011101100100011011011110000100110100110000;  // -2097447463 460868912
      11'h374: T=64'b1000001011110000101111011110100100011011010001110011001011101111;  // -2098151959 457650927
      11'h375: T=64'b1000001011100110000100010100001000011011000101100001010001111001;  // -2098851518 454431865
      11'h376: T=64'b1000001011011011011101111110011000011010111001001111000111010110;  // -2099546138 451211734
      11'h377: T=64'b1000001011010000111100011101011000011010101100111100101100001101;  // -2100235818 447990541
      11'h378: T=64'b1000001011000110011111110001010100011010100000101010000000100101;  // -2100920555 444768293
      11'h379: T=64'b1000001010111100000111111010001100011010010100010111000100101000;  // -2101600349 441545000
      11'h37a: T=64'b1000001010110001110100111000001000011010001000000011111000011011;  // -2102275198 438320667
      11'h37b: T=64'b1000001010100111100110101011010000011001111011110000011100000111;  // -2102945100 435095303
      11'h37c: T=64'b1000001010011101011101010011101100011001101111011100101111110011;  // -2103610053 431868915
      11'h37d: T=64'b1000001010010011011000110001100000011001100011001000110011100110;  // -2104270056 428641510
      11'h37e: T=64'b1000001010001001011001000100110000011001010110110100100111101010;  // -2104925108 425413098
      11'h37f: T=64'b1000001001111111011110001101100100011001001010100000001100000100;  // -2105575207 422183684
      11'h380: T=64'b1000001001110101101000001100000100011000111110001011100000111100;  // -2106220351 418953276
      11'h381: T=64'b1000001001101011110111000000010100011000110001110110100110011011;  // -2106860539 415721883
      11'h382: T=64'b1000001001100010001010101010011100011000100101100001011100101000;  // -2107495769 412489512
      11'h383: T=64'b1000001001011000100011001010100000011000011001001100000011101010;  // -2108126040 409256170
      11'h384: T=64'b1000001001001111000000100000100100011000001100110110011011101000;  // -2108751351 406021864
      11'h385: T=64'b1000001001000101100010101100110100011000000000100000100100101100;  // -2109371699 402786604
      11'h386: T=64'b1000001000111100001001101111010000010111110100001010011110111100;  // -2109987084 399550396
      11'h387: T=64'b1000001000110010110101101000000000010111100111110100001010011111;  // -2110597504 396313247
      11'h388: T=64'b1000001000101001100110010111001000010111011011011101100111011110;  // -2111202958 393075166
      11'h389: T=64'b1000001000100000011011111100110100010111001111000110110110000000;  // -2111803443 389836160
      11'h38a: T=64'b1000001000010111010110011001000100010111000010101111110110001101;  // -2112398959 386596237
      11'h38b: T=64'b1000001000001110010101101011111100010110110110011000101000001100;  // -2112989505 383355404
      11'h38c: T=64'b1000001000000101011001110101100100010110101010000001001100000101;  // -2113575079 380113669
      11'h38d: T=64'b1000000111111100100010110110000100010110011101101001100001111111;  // -2114155679 376871039
      11'h38e: T=64'b1000000111110011110000101101100000010110010001010001101010000011;  // -2114731304 373627523
      11'h38f: T=64'b1000000111101011000011011011111100010110000100111001100100010111;  // -2115301953 370383127
      11'h390: T=64'b1000000111100010011011000001011100010101111000100001010001000100;  // -2115867625 367137860
      11'h391: T=64'b1000000111011001110111011110001000010101101100001000110000010001;  // -2116428318 363891729
      11'h392: T=64'b1000000111010001011000110010001000010101011111110000000010000110;  // -2116984030 360644742
      11'h393: T=64'b1000000111001000111110111101011100010101010011010111000110101010;  // -2117534761 357396906
      11'h394: T=64'b1000000111000000101010000000001000010101000110111101111110000101;  // -2118080510 354148229
      11'h395: T=64'b1000000110111000011001111010011000010100111010100100101000011111;  // -2118621274 350898719
      11'h396: T=64'b1000000110110000001110101100001100010100101110001011000101111111;  // -2119157053 347648383
      11'h397: T=64'b1000000110101000001000010101101000010100100001110001010110101101;  // -2119687846 344397229
      11'h398: T=64'b1000000110100000000110110110111000010100010101010111011010110001;  // -2120213650 341145265
      11'h399: T=64'b1000000110011000001010001111111000010100001000111101010010010010;  // -2120734466 337892498
      11'h39a: T=64'b1000000110010000010010100000110100010011111100100010111101011000;  // -2121250291 334638936
      11'h39b: T=64'b1000000110001000011111101001101100010011110000001000011100001010;  // -2121761125 331384586
      11'h39c: T=64'b1000000110000000110001101010101000010011100011101101101110110001;  // -2122266966 328129457
      11'h39d: T=64'b1000000101111001001000100011101100010011010111010010110101010011;  // -2122767813 324873555
      11'h39e: T=64'b1000000101110001100100010100111100010011001010110111101111111001;  // -2123263665 321616889
      11'h39f: T=64'b1000000101101010000100111110011100010010111110011100011110101010;  // -2123754521 318359466
      11'h3a0: T=64'b1000000101100010101010100000010100010010110010000001000001101110;  // -2124240379 315101294
      11'h3a1: T=64'b1000000101011011010100111010100100010010100101100101011001001101;  // -2124721239 311842381
      11'h3a2: T=64'b1000000101010100000100001101010100010010011001001001100101001110;  // -2125197099 308582734
      11'h3a3: T=64'b1000000101001100111000011000100100010010001100101101100101111001;  // -2125667959 305322361
      11'h3a4: T=64'b1000000101000101110001011100100000010010000000010001011011010101;  // -2126133816 302061269
      11'h3a5: T=64'b1000000100111110101111011001000100010001110011110101000101101010;  // -2126594671 298799466
      11'h3a6: T=64'b1000000100110111110010001110011100010001100111011000100101000001;  // -2127050521 295536961
      11'h3a7: T=64'b1000000100110000111001111100101000010001011010111011111001100000;  // -2127501366 292273760
      11'h3a8: T=64'b1000000100101010000110100011101100010001001110011111000011001111;  // -2127947205 289009871
      11'h3a9: T=64'b1000000100100011011000000011101100010001000010000010000010010110;  // -2128388037 285745302
      11'h3aa: T=64'b1000000100011100101110011100101100010000110101100100110110111101;  // -2128823861 282480061
      11'h3ab: T=64'b1000000100010110001001101110110100010000101001000111100001001011;  // -2129254675 279214155
      11'h3ac: T=64'b1000000100001111101001111010000100010000011100101010000001001000;  // -2129680479 275947592
      11'h3ad: T=64'b1000000100001001001110111110100100010000010000001100010110111011;  // -2130101271 272680379
      11'h3ae: T=64'b1000000100000010111000111100010100010000000011101110100010101101;  // -2130517051 269412525
      11'h3af: T=64'b1000000011111100100111110011011000001111110111010000100100100101;  // -2130927818 266144037
      11'h3b0: T=64'b1000000011110110011011100011110100001111101010110010011100101011;  // -2131333571 262874923
      11'h3b1: T=64'b1000000011110000010100001101110000001111011110010100001011000110;  // -2131734308 259605190
      11'h3b2: T=64'b1000000011101010010001110001001100001111010001110101101111111111;  // -2132130029 256334847
      11'h3b3: T=64'b1000000011100100010100001110001100001111000101010111001011011100;  // -2132520733 253063900
      11'h3b4: T=64'b1000000011011110011011100100110100001110111000111000011101100110;  // -2132906419 249792358
      11'h3b5: T=64'b1000000011011000100111110101001000001110101100011001100110100100;  // -2133287086 246520228
      11'h3b6: T=64'b1000000011010010111000111111001100001110011111111010100110011101;  // -2133662733 243247517
      11'h3b7: T=64'b1000000011001101001111000011000000001110010011011011011101011011;  // -2134033360 239974235
      11'h3b8: T=64'b1000000011000111101010000000101100001110000110111100001011100100;  // -2134398965 236700388
      11'h3b9: T=64'b1000000011000010001001111000010100001101111010011100110000111111;  // -2134759547 233425983
      11'h3ba: T=64'b1000000010111100101110101001111000001101101101111101001101110110;  // -2135115106 230151030
      11'h3bb: T=64'b1000000010110111011000010101011100001101100001011101100010001111;  // -2135465641 226875535
      11'h3bc: T=64'b1000000010110010000110111011000000001101010100111101101110010010;  // -2135811152 223599506
      11'h3bd: T=64'b1000000010101100111010011010110000001101001000011101110010000111;  // -2136151636 220322951
      11'h3be: T=64'b1000000010100111110010110100101000001100111011111101101101110101;  // -2136487094 217045877
      11'h3bf: T=64'b1000000010100010110000001000110000001100101111011101100001100101;  // -2136817524 213768293
      11'h3c0: T=64'b1000000010011101110010010111001000001100100010111101001101011110;  // -2137142926 210490206
      11'h3c1: T=64'b1000000010011000111001011111110000001100010110011100110001100111;  // -2137463300 207211623
      11'h3c2: T=64'b1000000010010100000101100010110100001100001001111100001110001001;  // -2137778643 203932553
      11'h3c3: T=64'b1000000010001111010110100000001100001011111101011011100011001011;  // -2138088957 200653003
      11'h3c4: T=64'b1000000010001010101100011000000100001011110000111010110000110101;  // -2138394239 197372981
      11'h3c5: T=64'b1000000010000110000111001010011100001011100100011001110111001110;  // -2138694489 194092494
      11'h3c6: T=64'b1000000010000001100110110111010100001011010111111000110110011111;  // -2138989707 190811551
      11'h3c7: T=64'b1000000001111101001011011110110100001011001011010111101110101111;  // -2139279891 187530159
      11'h3c8: T=64'b1000000001111000110101000000111000001010111110110110100000000101;  // -2139565042 184248325
      11'h3c9: T=64'b1000000001110100100011011101101000001010110010010101001010101010;  // -2139845158 180966058
      11'h3ca: T=64'b1000000001110000010110110101000100001010100101110011101110100101;  // -2140120239 177683365
      11'h3cb: T=64'b1000000001101100001111000111010100001010011001010010001011111110;  // -2140390283 174400254
      11'h3cc: T=64'b1000000001101000001100010100010000001010001100110000100010111100;  // -2140655292 171116732
      11'h3cd: T=64'b1000000001100100001110011100000100001010000000001110110011101000;  // -2140915263 167832808
      11'h3ce: T=64'b1000000001100000010101011110110000001001110011101100111110001001;  // -2141170196 164548489
      11'h3cf: T=64'b1000000001011100100001011100010100001001100111001011000010100111;  // -2141420091 161263783
      11'h3d0: T=64'b1000000001011000110010010100110100001001011010101001000001001001;  // -2141664947 157978697
      11'h3d1: T=64'b1000000001010101001000001000010100001001001110000110111001111000;  // -2141904763 154693240
      11'h3d2: T=64'b1000000001010001100010110110110000001001000001100100101100111010;  // -2142139540 151407418
      11'h3d3: T=64'b1000000001001110000010100000010100001000110101000010011010011001;  // -2142369275 148121241
      11'h3d4: T=64'b1000000001001010100111000100111000001000101000100000000010011010;  // -2142593970 144834714
      11'h3d5: T=64'b1000000001000111010000100100100100001000011011111101100101000111;  // -2142813623 141547847
      11'h3d6: T=64'b1000000001000011111110111111011100001000001111011011000010100111;  // -2143028233 138260647
      11'h3d7: T=64'b1000000001000000110010010101011100001000000010111000011011000010;  // -2143237801 134973122
      11'h3d8: T=64'b1000000000111101101010100110101100000111110110010101101110011110;  // -2143442325 131685278
      11'h3d9: T=64'b1000000000111010100111110011001000000111101001110010111101000101;  // -2143641806 128397125
      11'h3da: T=64'b1000000000110111101001111010110100000111011101010000000110111110;  // -2143836243 125108670
      11'h3db: T=64'b1000000000110100110000111101111000000111010000101101001100010001;  // -2144025634 121819921
      11'h3dc: T=64'b1000000000110001111100111100001100000111000100001010001101000101;  // -2144209981 118530885
      11'h3dd: T=64'b1000000000101111001101110101111000000110110111100111001001100010;  // -2144389282 115241570
      11'h3de: T=64'b1000000000101100100011101010111000000110101011000100000001101111;  // -2144563538 111951983
      11'h3df: T=64'b1000000000101001111110011011010100000110011110100000110101110110;  // -2144732747 108662134
      11'h3e0: T=64'b1000000000100111011110000111001100000110010001111101100101111100;  // -2144896909 105372028
      11'h3e1: T=64'b1000000000100101000010101110100000000110000101011010010010001011;  // -2145056024 102081675
      11'h3e2: T=64'b1000000000100010101100010001010100000101111000110110111010101001;  // -2145210091 98791081
      11'h3e3: T=64'b1000000000100000011010101111100100000101101100010011011111011111;  // -2145359111 95500255
      11'h3e4: T=64'b1000000000011110001110001001011000000101011111110000000000110101;  // -2145503082 92209205
      11'h3e5: T=64'b1000000000011100000110011110101100000101010011001100011110110001;  // -2145642005 88917937
      11'h3e6: T=64'b1000000000011010000011101111100100000101000110101000111001011100;  // -2145775879 85626460
      11'h3e7: T=64'b1000000000011000000101111100000000000100111010000101010000111110;  // -2145904704 82334782
      11'h3e8: T=64'b1000000000010110001101000100000100000100101101100001100101011101;  // -2146028479 79042909
      11'h3e9: T=64'b1000000000010100011001000111110000000100100000111101110111000011;  // -2146147204 75750851
      11'h3ea: T=64'b1000000000010010101010000111000000000100010100011010000101110111;  // -2146260880 72458615
      11'h3eb: T=64'b1000000000010001000000000010000000000100000111110110010010000000;  // -2146369504 69166208
      11'h3ec: T=64'b1000000000001111011010111000100100000011111011010010011011100110;  // -2146473079 65873638
      11'h3ed: T=64'b1000000000001101111010101010111000000011101110101110100010110010;  // -2146571602 62580914
      11'h3ee: T=64'b1000000000001100011111011000110100000011100010001010100111101010;  // -2146665075 59288042
      11'h3ef: T=64'b1000000000001011001001000010100000000011010101100110101010010110;  // -2146753496 55995030
      11'h3f0: T=64'b1000000000001001110111100111111100000011001001000010101010111111;  // -2146836865 52701887
      11'h3f1: T=64'b1000000000001000101011001001000100000010111100011110101001101100;  // -2146915183 49408620
      11'h3f2: T=64'b1000000000000111100011100101111100000010101111111010100110100100;  // -2146988449 46115236
      11'h3f3: T=64'b1000000000000110100000111110100100000010100011010110100001110000;  // -2147056663 42821744
      11'h3f4: T=64'b1000000000000101100011010011000000000010010110110010011011010111;  // -2147119824 39528151
      11'h3f5: T=64'b1000000000000100101010100011001100000010001010001110010011100010;  // -2147177933 36234466
      11'h3f6: T=64'b1000000000000011110110101111001000000001111101101010001010010111;  // -2147230990 32940695
      11'h3f7: T=64'b1000000000000011000111110110111000000001110001000101111111111110;  // -2147278994 29646846
      11'h3f8: T=64'b1000000000000010011101111010011100000001100100100001110100100000;  // -2147321945 26352928
      11'h3f9: T=64'b1000000000000001111000111001110000000001010111111101101000000011;  // -2147359844 23058947
      11'h3fa: T=64'b1000000000000001011000110100111100000001001011011001011010110001;  // -2147392689 19764913
      11'h3fb: T=64'b1000000000000000111101101011111000000000111110110101001100110000;  // -2147420482 16470832
      11'h3fc: T=64'b1000000000000000100111011110101100000000110010010000111110001000;  // -2147443221 13176712
      11'h3fd: T=64'b1000000000000000010110001101010100000000100101101100101111000001;  // -2147460907 9882561
      11'h3fe: T=64'b1000000000000000001001110111101100000000011001001000011111100011;  // -2147473541 6588387
      11'h3ff: T=64'b1000000000000000000010011110000000000000001100100100001111110101;  // -2147481120 3294197
      11'h400: T=64'b1000000000000000000000000000000100000000000000000000000000000000;  // -2147483647     0
      11'h401: T=64'b1000000000000000000010011110000011111111110011011011110000001011;  // -2147481120 -3294197
      11'h402: T=64'b1000000000000000001001110111101111111111100110110111100000011101;  // -2147473541 -6588387
      11'h403: T=64'b1000000000000000010110001101010111111111011010010011010000111111;  // -2147460907 -9882561
      11'h404: T=64'b1000000000000000100111011110101111111111001101101111000001111000;  // -2147443221 -13176712
      11'h405: T=64'b1000000000000000111101101011111011111111000001001010110011010000;  // -2147420482 -16470832
      11'h406: T=64'b1000000000000001011000110100111111111110110100100110100101001111;  // -2147392689 -19764913
      11'h407: T=64'b1000000000000001111000111001110011111110101000000010010111111101;  // -2147359844 -23058947
      11'h408: T=64'b1000000000000010011101111010011111111110011011011110001011100000;  // -2147321945 -26352928
      11'h409: T=64'b1000000000000011000111110110111011111110001110111010000000000010;  // -2147278994 -29646846
      11'h40a: T=64'b1000000000000011110110101111001011111110000010010101110101101001;  // -2147230990 -32940695
      11'h40b: T=64'b1000000000000100101010100011001111111101110101110001101100011110;  // -2147177933 -36234466
      11'h40c: T=64'b1000000000000101100011010011000011111101101001001101100100101001;  // -2147119824 -39528151
      11'h40d: T=64'b1000000000000110100000111110100111111101011100101001011110010000;  // -2147056663 -42821744
      11'h40e: T=64'b1000000000000111100011100101111111111101010000000101011001011100;  // -2146988449 -46115236
      11'h40f: T=64'b1000000000001000101011001001000111111101000011100001010110010100;  // -2146915183 -49408620
      11'h410: T=64'b1000000000001001110111100111111111111100110110111101010101000001;  // -2146836865 -52701887
      11'h411: T=64'b1000000000001011001001000010100011111100101010011001010101101010;  // -2146753496 -55995030
      11'h412: T=64'b1000000000001100011111011000110111111100011101110101011000010110;  // -2146665075 -59288042
      11'h413: T=64'b1000000000001101111010101010111011111100010001010001011101001110;  // -2146571602 -62580914
      11'h414: T=64'b1000000000001111011010111000100111111100000100101101100100011010;  // -2146473079 -65873638
      11'h415: T=64'b1000000000010001000000000010000011111011111000001001101110000000;  // -2146369504 -69166208
      11'h416: T=64'b1000000000010010101010000111000011111011101011100101111010001001;  // -2146260880 -72458615
      11'h417: T=64'b1000000000010100011001000111110011111011011111000010001000111101;  // -2146147204 -75750851
      11'h418: T=64'b1000000000010110001101000100000111111011010010011110011010100011;  // -2146028479 -79042909
      11'h419: T=64'b1000000000011000000101111100000011111011000101111010101111000010;  // -2145904704 -82334782
      11'h41a: T=64'b1000000000011010000011101111100111111010111001010111000110100100;  // -2145775879 -85626460
      11'h41b: T=64'b1000000000011100000110011110101111111010101100110011100001001111;  // -2145642005 -88917937
      11'h41c: T=64'b1000000000011110001110001001011011111010100000001111111111001011;  // -2145503082 -92209205
      11'h41d: T=64'b1000000000100000011010101111100111111010010011101100100000100001;  // -2145359111 -95500255
      11'h41e: T=64'b1000000000100010101100010001010111111010000111001001000101010111;  // -2145210091 -98791081
      11'h41f: T=64'b1000000000100101000010101110100011111001111010100101101101110101;  // -2145056024 -102081675
      11'h420: T=64'b1000000000100111011110000111001111111001101110000010011010000100;  // -2144896909 -105372028
      11'h421: T=64'b1000000000101001111110011011010111111001100001011111001010001010;  // -2144732747 -108662134
      11'h422: T=64'b1000000000101100100011101010111011111001010100111011111110010001;  // -2144563538 -111951983
      11'h423: T=64'b1000000000101111001101110101111011111001001000011000110110011110;  // -2144389282 -115241570
      11'h424: T=64'b1000000000110001111100111100001111111000111011110101110010111011;  // -2144209981 -118530885
      11'h425: T=64'b1000000000110100110000111101111011111000101111010010110011101111;  // -2144025634 -121819921
      11'h426: T=64'b1000000000110111101001111010110111111000100010101111111001000010;  // -2143836243 -125108670
      11'h427: T=64'b1000000000111010100111110011001011111000010110001101000010111011;  // -2143641806 -128397125
      11'h428: T=64'b1000000000111101101010100110101111111000001001101010010001100010;  // -2143442325 -131685278
      11'h429: T=64'b1000000001000000110010010101011111110111111101000111100100111110;  // -2143237801 -134973122
      11'h42a: T=64'b1000000001000011111110111111011111110111110000100100111101011001;  // -2143028233 -138260647
      11'h42b: T=64'b1000000001000111010000100100100111110111100100000010011010111001;  // -2142813623 -141547847
      11'h42c: T=64'b1000000001001010100111000100111011110111010111011111111101100110;  // -2142593970 -144834714
      11'h42d: T=64'b1000000001001110000010100000010111110111001010111101100101100111;  // -2142369275 -148121241
      11'h42e: T=64'b1000000001010001100010110110110011110110111110011011010011000110;  // -2142139540 -151407418
      11'h42f: T=64'b1000000001010101001000001000010111110110110001111001000110001000;  // -2141904763 -154693240
      11'h430: T=64'b1000000001011000110010010100110111110110100101010110111110110111;  // -2141664947 -157978697
      11'h431: T=64'b1000000001011100100001011100010111110110011000110100111101011001;  // -2141420091 -161263783
      11'h432: T=64'b1000000001100000010101011110110011110110001100010011000001110111;  // -2141170196 -164548489
      11'h433: T=64'b1000000001100100001110011100000111110101111111110001001100011000;  // -2140915263 -167832808
      11'h434: T=64'b1000000001101000001100010100010011110101110011001111011101000100;  // -2140655292 -171116732
      11'h435: T=64'b1000000001101100001111000111010111110101100110101101110100000010;  // -2140390283 -174400254
      11'h436: T=64'b1000000001110000010110110101000111110101011010001100010001011011;  // -2140120239 -177683365
      11'h437: T=64'b1000000001110100100011011101101011110101001101101010110101010110;  // -2139845158 -180966058
      11'h438: T=64'b1000000001111000110101000000111011110101000001001001011111111011;  // -2139565042 -184248325
      11'h439: T=64'b1000000001111101001011011110110111110100110100101000010001010001;  // -2139279891 -187530159
      11'h43a: T=64'b1000000010000001100110110111010111110100101000000111001001100001;  // -2138989707 -190811551
      11'h43b: T=64'b1000000010000110000111001010011111110100011011100110001000110010;  // -2138694489 -194092494
      11'h43c: T=64'b1000000010001010101100011000000111110100001111000101001111001011;  // -2138394239 -197372981
      11'h43d: T=64'b1000000010001111010110100000001111110100000010100100011100110101;  // -2138088957 -200653003
      11'h43e: T=64'b1000000010010100000101100010110111110011110110000011110001110111;  // -2137778643 -203932553
      11'h43f: T=64'b1000000010011000111001011111110011110011101001100011001110011001;  // -2137463300 -207211623
      11'h440: T=64'b1000000010011101110010010111001011110011011101000010110010100010;  // -2137142926 -210490206
      11'h441: T=64'b1000000010100010110000001000110011110011010000100010011110011011;  // -2136817524 -213768293
      11'h442: T=64'b1000000010100111110010110100101011110011000100000010010010001011;  // -2136487094 -217045877
      11'h443: T=64'b1000000010101100111010011010110011110010110111100010001101111001;  // -2136151636 -220322951
      11'h444: T=64'b1000000010110010000110111011000011110010101011000010010001101110;  // -2135811152 -223599506
      11'h445: T=64'b1000000010110111011000010101011111110010011110100010011101110001;  // -2135465641 -226875535
      11'h446: T=64'b1000000010111100101110101001111011110010010010000010110010001010;  // -2135115106 -230151030
      11'h447: T=64'b1000000011000010001001111000010111110010000101100011001111000001;  // -2134759547 -233425983
      11'h448: T=64'b1000000011000111101010000000101111110001111001000011110100011100;  // -2134398965 -236700388
      11'h449: T=64'b1000000011001101001111000011000011110001101100100100100010100101;  // -2134033360 -239974235
      11'h44a: T=64'b1000000011010010111000111111001111110001100000000101011001100011;  // -2133662733 -243247517
      11'h44b: T=64'b1000000011011000100111110101001011110001010011100110011001011100;  // -2133287086 -246520228
      11'h44c: T=64'b1000000011011110011011100100110111110001000111000111100010011010;  // -2132906419 -249792358
      11'h44d: T=64'b1000000011100100010100001110001111110000111010101000110100100100;  // -2132520733 -253063900
      11'h44e: T=64'b1000000011101010010001110001001111110000101110001010010000000001;  // -2132130029 -256334847
      11'h44f: T=64'b1000000011110000010100001101110011110000100001101011110100111010;  // -2131734308 -259605190
      11'h450: T=64'b1000000011110110011011100011110111110000010101001101100011010101;  // -2131333571 -262874923
      11'h451: T=64'b1000000011111100100111110011011011110000001000101111011011011011;  // -2130927818 -266144037
      11'h452: T=64'b1000000100000010111000111100010111101111111100010001011101010011;  // -2130517051 -269412525
      11'h453: T=64'b1000000100001001001110111110100111101111101111110011101001000101;  // -2130101271 -272680379
      11'h454: T=64'b1000000100001111101001111010000111101111100011010101111110111000;  // -2129680479 -275947592
      11'h455: T=64'b1000000100010110001001101110110111101111010110111000011110110101;  // -2129254675 -279214155
      11'h456: T=64'b1000000100011100101110011100101111101111001010011011001001000011;  // -2128823861 -282480061
      11'h457: T=64'b1000000100100011011000000011101111101110111101111101111101101010;  // -2128388037 -285745302
      11'h458: T=64'b1000000100101010000110100011101111101110110001100000111100110001;  // -2127947205 -289009871
      11'h459: T=64'b1000000100110000111001111100101011101110100101000100000110100000;  // -2127501366 -292273760
      11'h45a: T=64'b1000000100110111110010001110011111101110011000100111011010111111;  // -2127050521 -295536961
      11'h45b: T=64'b1000000100111110101111011001000111101110001100001010111010010110;  // -2126594671 -298799466
      11'h45c: T=64'b1000000101000101110001011100100011101101111111101110100100101011;  // -2126133816 -302061269
      11'h45d: T=64'b1000000101001100111000011000100111101101110011010010011010000111;  // -2125667959 -305322361
      11'h45e: T=64'b1000000101010100000100001101010111101101100110110110011010110010;  // -2125197099 -308582734
      11'h45f: T=64'b1000000101011011010100111010100111101101011010011010100110110011;  // -2124721239 -311842381
      11'h460: T=64'b1000000101100010101010100000010111101101001101111110111110010010;  // -2124240379 -315101294
      11'h461: T=64'b1000000101101010000100111110011111101101000001100011100001010110;  // -2123754521 -318359466
      11'h462: T=64'b1000000101110001100100010100111111101100110101001000010000000111;  // -2123263665 -321616889
      11'h463: T=64'b1000000101111001001000100011101111101100101000101101001010101101;  // -2122767813 -324873555
      11'h464: T=64'b1000000110000000110001101010101011101100011100010010010001001111;  // -2122266966 -328129457
      11'h465: T=64'b1000000110001000011111101001101111101100001111110111100011110110;  // -2121761125 -331384586
      11'h466: T=64'b1000000110010000010010100000110111101100000011011101000010101000;  // -2121250291 -334638936
      11'h467: T=64'b1000000110011000001010001111111011101011110111000010101101101110;  // -2120734466 -337892498
      11'h468: T=64'b1000000110100000000110110110111011101011101010101000100101001111;  // -2120213650 -341145265
      11'h469: T=64'b1000000110101000001000010101101011101011011110001110101001010011;  // -2119687846 -344397229
      11'h46a: T=64'b1000000110110000001110101100001111101011010001110100111010000001;  // -2119157053 -347648383
      11'h46b: T=64'b1000000110111000011001111010011011101011000101011011010111100001;  // -2118621274 -350898719
      11'h46c: T=64'b1000000111000000101010000000001011101010111001000010000001111011;  // -2118080510 -354148229
      11'h46d: T=64'b1000000111001000111110111101011111101010101100101000111001010110;  // -2117534761 -357396906
      11'h46e: T=64'b1000000111010001011000110010001011101010100000001111111101111010;  // -2116984030 -360644742
      11'h46f: T=64'b1000000111011001110111011110001011101010010011110111001111101111;  // -2116428318 -363891729
      11'h470: T=64'b1000000111100010011011000001011111101010000111011110101110111100;  // -2115867625 -367137860
      11'h471: T=64'b1000000111101011000011011011111111101001111011000110011011101001;  // -2115301953 -370383127
      11'h472: T=64'b1000000111110011110000101101100011101001101110101110010101111101;  // -2114731304 -373627523
      11'h473: T=64'b1000000111111100100010110110000111101001100010010110011110000001;  // -2114155679 -376871039
      11'h474: T=64'b1000001000000101011001110101100111101001010101111110110011111011;  // -2113575079 -380113669
      11'h475: T=64'b1000001000001110010101101011111111101001001001100111010111110100;  // -2112989505 -383355404
      11'h476: T=64'b1000001000010111010110011001000111101000111101010000001001110011;  // -2112398959 -386596237
      11'h477: T=64'b1000001000100000011011111100110111101000110000111001001010000000;  // -2111803443 -389836160
      11'h478: T=64'b1000001000101001100110010111001011101000100100100010011000100010;  // -2111202958 -393075166
      11'h479: T=64'b1000001000110010110101101000000011101000011000001011110101100001;  // -2110597504 -396313247
      11'h47a: T=64'b1000001000111100001001101111010011101000001011110101100001000100;  // -2109987084 -399550396
      11'h47b: T=64'b1000001001000101100010101100110111100111111111011111011011010100;  // -2109371699 -402786604
      11'h47c: T=64'b1000001001001111000000100000100111100111110011001001100100011000;  // -2108751351 -406021864
      11'h47d: T=64'b1000001001011000100011001010100011100111100110110011111100010110;  // -2108126040 -409256170
      11'h47e: T=64'b1000001001100010001010101010011111100111011010011110100011011000;  // -2107495769 -412489512
      11'h47f: T=64'b1000001001101011110111000000010111100111001110001001011001100101;  // -2106860539 -415721883
      11'h480: T=64'b1000001001110101101000001100000111100111000001110100011111000100;  // -2106220351 -418953276
      11'h481: T=64'b1000001001111111011110001101100111100110110101011111110011111100;  // -2105575207 -422183684
      11'h482: T=64'b1000001010001001011001000100110011100110101001001011011000010110;  // -2104925108 -425413098
      11'h483: T=64'b1000001010010011011000110001100011100110011100110111001100011010;  // -2104270056 -428641510
      11'h484: T=64'b1000001010011101011101010011101111100110010000100011010000001101;  // -2103610053 -431868915
      11'h485: T=64'b1000001010100111100110101011010011100110000100001111100011111001;  // -2102945100 -435095303
      11'h486: T=64'b1000001010110001110100111000001011100101110111111100000111100101;  // -2102275198 -438320667
      11'h487: T=64'b1000001010111100000111111010001111100101101011101000111011011000;  // -2101600349 -441545000
      11'h488: T=64'b1000001011000110011111110001010111100101011111010101111111011011;  // -2100920555 -444768293
      11'h489: T=64'b1000001011010000111100011101011011100101010011000011010011110011;  // -2100235818 -447990541
      11'h48a: T=64'b1000001011011011011101111110011011100101000110110000111000101010;  // -2099546138 -451211734
      11'h48b: T=64'b1000001011100110000100010100001011100100111010011110101110000111;  // -2098851518 -454431865
      11'h48c: T=64'b1000001011110000101111011110100111100100101110001100110100010001;  // -2098151959 -457650927
      11'h48d: T=64'b1000001011111011011111011101100111100100100001111011001011010000;  // -2097447463 -460868912
      11'h48e: T=64'b1000001100000110010100010001000111100100010101101001110011001011;  // -2096738031 -464085813
      11'h48f: T=64'b1000001100010001001101111000111011100100001001011000101100001011;  // -2096023666 -467301621
      11'h490: T=64'b1000001100011100001100010100111111100011111101000111110110010110;  // -2095304369 -470516330
      11'h491: T=64'b1000001100100111001111100101001111100011110000110111010001110100;  // -2094580141 -473729932
      11'h492: T=64'b1000001100110010010111101001100011100011100100100110111110101101;  // -2093850984 -476942419
      11'h493: T=64'b1000001100111101100100100001110011100011011000010110111101001000;  // -2093116900 -480153784
      11'h494: T=64'b1000001101001000110110001101110111100011001100000111001101001101;  // -2092377891 -483364019
      11'h495: T=64'b1000001101010100001100101101100111100010111111110111101111000100;  // -2091633959 -486573116
      11'h496: T=64'b1000001101011111101000000001000011100010110011101000100010110011;  // -2090885104 -489781069
      11'h497: T=64'b1000001101101011001000000111111011100010100111011001101000100011;  // -2090131330 -492987869
      11'h498: T=64'b1000001101110110101101000010001111100010011011001011000000011011;  // -2089372637 -496193509
      11'h499: T=64'b1000001110000010010110101111110011100010001110111100101010100011;  // -2088609028 -499397981
      11'h49a: T=64'b1000001110001110000101010000100011100010000010101110100111000001;  // -2087840504 -502601279
      11'h49b: T=64'b1000001110011001111000100100010111100001110110100000110101111111;  // -2087067067 -505803393
      11'h49c: T=64'b1000001110100101110000101011000111100001101010010011010111100010;  // -2086288719 -509004318
      11'h49d: T=64'b1000001110110001101101100100101011100001011110000110001011110011;  // -2085505462 -512204045
      11'h49e: T=64'b1000001110111101101111010000111111100001010001111001010010111010;  // -2084717297 -515402566
      11'h49f: T=64'b1000001111001001110101101111110111100001000101101100101100111101;  // -2083924227 -518599875
      11'h4a0: T=64'b1000001111010110000001000001001111100000111001100000011010000101;  // -2083126253 -521795963
      11'h4a1: T=64'b1000001111100010010001000100111011100000101101010100011010011001;  // -2082323378 -524990823
      11'h4a2: T=64'b1000001111101110100101111010111011100000100001001000101110000000;  // -2081515602 -528184448
      11'h4a3: T=64'b1000001111111010111111100010111111100000010100111101010101000001;  // -2080702929 -531376831
      11'h4a4: T=64'b1000010000000111011101111101000111100000001000110010001111100101;  // -2079885359 -534567963
      11'h4a5: T=64'b1000010000010100000001001001000111011111111100100111011101110011;  // -2079062895 -537757837
      11'h4a6: T=64'b1000010000100000101001000110110111011111110000011100111111110011;  // -2078235539 -540946445
      11'h4a7: T=64'b1000010000101101010101110110001111011111100100010010110101101011;  // -2077403293 -544133781
      11'h4a8: T=64'b1000010000111010000111010111000111011111011000001000111111100100;  // -2076566159 -547319836
      11'h4a9: T=64'b1000010001000110111101101001011011011111001011111111011101100100;  // -2075724138 -550504604
      11'h4aa: T=64'b1000010001010011111000101101000011011110111111110110001111110100;  // -2074877232 -553688076
      11'h4ab: T=64'b1000010001100000111000100001101111011110110011101101010110011011;  // -2074025445 -556870245
      11'h4ac: T=64'b1000010001101101111101000111100011011110100111100100110001100001;  // -2073168776 -560051103
      11'h4ad: T=64'b1000010001111011000110011110001011011110011011011100100001001100;  // -2072307230 -563230644
      11'h4ae: T=64'b1000010010001000010100100101100111011110001111010100100101100100;  // -2071440807 -566408860
      11'h4af: T=64'b1000010010010101100111011101101011011110000011001100111110110001;  // -2070569510 -569585743
      11'h4b0: T=64'b1000010010100010111111000110001111011101110111000101101100111011;  // -2069693341 -572761285
      11'h4b1: T=64'b1000010010110000011011011111001111011101101010111110110000001000;  // -2068812301 -575935480
      11'h4b2: T=64'b1000010010111101111100101000011111011101011110111000001000100001;  // -2067926393 -579108319
      11'h4b3: T=64'b1000010011001011100010100001110011011101010010110001110110001100;  // -2067035620 -582279796
      11'h4b4: T=64'b1000010011011001001101001011001011011101000110101011111001010001;  // -2066139982 -585449903
      11'h4b5: T=64'b1000010011100110111100100100010111011100111010100110010001111000;  // -2065239483 -588618632
      11'h4b6: T=64'b1000010011110100110000101101010111011100101110100001000000001000;  // -2064334123 -591785976
      11'h4b7: T=64'b1000010100000010101001100101110111011100100010011100000100001001;  // -2063423907 -594951927
      11'h4b8: T=64'b1000010100010000100111001101110111011100010110010111011110000010;  // -2062508835 -598116478
      11'h4b9: T=64'b1000010100011110101001100101001111011100001010010011001101111010;  // -2061588909 -601279622
      11'h4ba: T=64'b1000010100101100110000101011110011011011111110001111010011111001;  // -2060664132 -604441351
      11'h4bb: T=64'b1000010100111010111100100001010111011011110010001011110000000110;  // -2059734507 -607601658
      11'h4bc: T=64'b1000010101001001001101000101110111011011100110001000100010101001;  // -2058800035 -610760535
      11'h4bd: T=64'b1000010101010111100010011001001011011011011010000101101011101001;  // -2057860718 -613917975
      11'h4be: T=64'b1000010101100101111100011011000111011011001110000011001011001110;  // -2056916559 -617073970
      11'h4bf: T=64'b1000010101110100011011001011100111011011000010000001000001011110;  // -2055967559 -620228514
      11'h4c0: T=64'b1000010110000010111110101010011011011010110101111111001110100011;  // -2055013722 -623381597
      11'h4c1: T=64'b1000010110010001100110110111011111011010101001111101110010100010;  // -2054055049 -626533214
      11'h4c2: T=64'b1000010110100000010011110010100111011010011101111100101101100011;  // -2053091543 -629683357
      11'h4c3: T=64'b1000010110101111000101011011101011011010010001111011111111101110;  // -2052123206 -632832018
      11'h4c4: T=64'b1000010110111101111011110010100011011010000101111011101001001010;  // -2051150040 -635979190
      11'h4c5: T=64'b1000010111001100110110110111000111011001111001111011101001111111;  // -2050172047 -639124865
      11'h4c6: T=64'b1000010111011011110110101001001011011001101101111100000010010100;  // -2049189230 -642269036
      11'h4c7: T=64'b1000010111101010111011001000100111011001100001111100110010010000;  // -2048201591 -645411696
      11'h4c8: T=64'b1000010111111010000100010101010011011001010101111101111001111011;  // -2047209132 -648552837
      11'h4c9: T=64'b1000011000001001010010001111000011011001001001111111011001011011;  // -2046211856 -651692453
      11'h4ca: T=64'b1000011000011000100100110101101011011000111110000001010000111010;  // -2045209766 -654830534
      11'h4cb: T=64'b1000011000100111111100001001001011011000110010000011100000011101;  // -2044202862 -657967075
      11'h4cc: T=64'b1000011000110111011000001001001111011000100110000110001000001100;  // -2043191149 -661102068
      11'h4cd: T=64'b1000011001000110111000110101110111011000011010001001001000001111;  // -2042174627 -664235505
      11'h4ce: T=64'b1000011001010110011110001110101111011000001110001100100000101101;  // -2041153301 -667367379
      11'h4cf: T=64'b1000011001100110001000010011110111011000000010010000010001101110;  // -2040127171 -670497682
      11'h4d0: T=64'b1000011001110101110111000101000011010111110110010100011011011000;  // -2039096240 -673626408
      11'h4d1: T=64'b1000011010000101101010100010000011010111101010011000111101110011;  // -2038060512 -676753549
      11'h4d2: T=64'b1000011010010101100010101010110111010111011110011101111001000111;  // -2037019987 -679879097
      11'h4d3: T=64'b1000011010100101011111011111001111010111010010100011001101011011;  // -2035974669 -683003045
      11'h4d4: T=64'b1000011010110101100000111110111111010111000110101000111010110110;  // -2034924561 -686125386
      11'h4d5: T=64'b1000011011000101100111001010000011010110111010101111000001011111;  // -2033869664 -689246113
      11'h4d6: T=64'b1000011011010101110010000000001111010110101110110101100001011110;  // -2032809981 -692365218
      11'h4d7: T=64'b1000011011100110000001100001010111010110100010111100011010111010;  // -2031745515 -695482694
      11'h4d8: T=64'b1000011011110110010101101101010011010110010111000011101101111011;  // -2030676268 -698598533
      11'h4d9: T=64'b1000011100000110101110100011111011010110001011001011011010101000;  // -2029602242 -701712728
      11'h4da: T=64'b1000011100010111001100000100111111010101111111010011100001001000;  // -2028523441 -704825272
      11'h4db: T=64'b1000011100100111101110010000011011010101110011011100000001100011;  // -2027439866 -707936157
      11'h4dc: T=64'b1000011100111000010101000101111111010101100111100100111011111111;  // -2026351521 -711045377
      11'h4dd: T=64'b1000011101001001000000100101100111010101011011101110010000100100;  // -2025258407 -714152924
      11'h4de: T=64'b1000011101011001110000101111000011010101001111110111111111011010;  // -2024160528 -717258790
      11'h4df: T=64'b1000011101101010100101100010001011010101000100000010001000101000;  // -2023057886 -720362968
      11'h4e0: T=64'b1000011101111011011110111110110111010100111000001100101100010101;  // -2021950483 -723465451
      11'h4e1: T=64'b1000011110001100011101000100111011010100101100010111101010101000;  // -2020838322 -726566232
      11'h4e2: T=64'b1000011110011101011111110100000111010100100000100011000011101001;  // -2019721407 -729665303
      11'h4e3: T=64'b1000011110101110100111001100011011010100010100101110110111011111;  // -2018599738 -732762657
      11'h4e4: T=64'b1000011110111111110011001101100011010100001000111011000110010001;  // -2017473320 -735858287
      11'h4e5: T=64'b1000011111010001000011110111011011010011111101000111110000000111;  // -2016342154 -738952185
      11'h4e6: T=64'b1000011111100010011001001001110011010011110001010100110101000111;  // -2015206244 -742044345
      11'h4e7: T=64'b1000011111110011110011000100100111010011100101100010010101011010;  // -2014065591 -745134758
      11'h4e8: T=64'b1000100000000101010001100111100011010011011001110000010001000110;  // -2012920200 -748223418
      11'h4e9: T=64'b1000100000010110110100110010100011010011001101111110101000010010;  // -2011770072 -751310318
      11'h4ea: T=64'b1000100000101000011100100101011111010011000010001101011011000111;  // -2010615209 -754395449
      11'h4eb: T=64'b1000100000111010001001000000000011010010110110011100101001101011;  // -2009455616 -757478805
      11'h4ec: T=64'b1000100001001011111010000010000111010010101010101100010100000101;  // -2008291295 -760560379
      11'h4ed: T=64'b1000100001011101101111101011100111010010011110111100011010011101;  // -2007122247 -763640163
      11'h4ee: T=64'b1000100001101111101001111100001111010010010011001100111100111001;  // -2005948477 -766718151
      11'h4ef: T=64'b1000100010000001101000110011111011010010000111011101111011100010;  // -2004769986 -769794334
      11'h4f0: T=64'b1000100010010011101100010010011011010001111011101111010110011110;  // -2003586778 -772868706
      11'h4f1: T=64'b1000100010100101110100010111100011010001110000000001001101110101;  // -2002398856 -775941259
      11'h4f2: T=64'b1000100010111000000001000011001111010001100100010011100001101110;  // -2001206221 -779011986
      11'h4f3: T=64'b1000100011001010010010010101001011010001011000100110010010010000;  // -2000008878 -782080880
      11'h4f4: T=64'b1000100011011100101000001101010011010001001100111001011111100010;  // -1998806828 -785147934
      11'h4f5: T=64'b1000100011101111000010101011010111010001000001001101001001101100;  // -1997600075 -788213140
      11'h4f6: T=64'b1000100100000001100001101111001111010000110101100001010000110100;  // -1996388621 -791276492
      11'h4f7: T=64'b1000100100010100000101011000101011010000101001110101110101000011;  // -1995172470 -794337981
      11'h4f8: T=64'b1000100100100110101101100111100011010000011110001010110110011110;  // -1993951624 -797397602
      11'h4f9: T=64'b1000100100111001011010011011101011010000010010100000010101001110;  // -1992726086 -800455346
      11'h4fa: T=64'b1000100101001100001011110100110111010000000110110110010001011001;  // -1991495859 -803511207
      11'h4fb: T=64'b1000100101011111000001110010111111001111111011001100101011001000;  // -1990260945 -806565176
      11'h4fc: T=64'b1000100101110001111100010101101111001111101111100011100010100000;  // -1989021349 -809617248
      11'h4fd: T=64'b1000100110000100111011011101000011001111100011111010110111101001;  // -1987777072 -812667415
      11'h4fe: T=64'b1000100110010111111111001000101111001111011000010010101010101010;  // -1986528117 -815715670
      11'h4ff: T=64'b1000100110101011000111011000100011001111001100101010111011101011;  // -1985274488 -818762005
      11'h500: T=64'b1000100110111110010100001100010011001111000001000011101010110011;  // -1984016188 -821806413
      11'h501: T=64'b1000100111010001100101100011110111001110110101011100111000001000;  // -1982753219 -824848888
      11'h502: T=64'b1000100111100100111011011111000011001110101001110110100011110011;  // -1981485584 -827889421
      11'h503: T=64'b1000100111111000010101111101100111001110011110010000101101111001;  // -1980213287 -830928007
      11'h504: T=64'b1000101000001011110100111111011011001110010010101011010110100011;  // -1978936330 -833964637
      11'h505: T=64'b1000101000011111011000100100010011001110000111000110011101110111;  // -1977654716 -836999305
      11'h506: T=64'b1000101000110011000000101011111111001101111011100010000011111101;  // -1976368449 -840032003
      11'h507: T=64'b1000101001000110101101010110010011001101101111111110001000111011;  // -1975077532 -843062725
      11'h508: T=64'b1000101001011010011110100011001011001101100100011010101100111001;  // -1973781966 -846091463
      11'h509: T=64'b1000101001101110010100010010010011001101011000110111101111111110;  // -1972481756 -849118210
      11'h50a: T=64'b1000101010000010001110100011011111001101001101010101010010010001;  // -1971176905 -852142959
      11'h50b: T=64'b1000101010010110001101010110100011001101000001110011010011111001;  // -1969867416 -855165703
      11'h50c: T=64'b1000101010101010010000101011010111001100110110010001110100111110;  // -1968553291 -858186434
      11'h50d: T=64'b1000101010111110011000100001101011001100101010110000110101100110;  // -1967234534 -861205146
      11'h50e: T=64'b1000101011010010100100111001010111001100011111010000010101111000;  // -1965911147 -864221832
      11'h50f: T=64'b1000101011100110110101110010000111001100010011110000010101111100;  // -1964583135 -867236484
      11'h510: T=64'b1000101011111011001011001011110011001100001000010000110101111001;  // -1963250500 -870249095
      11'h511: T=64'b1000101100001111100101000110001011001011111100110001110101110110;  // -1961913246 -873259658
      11'h512: T=64'b1000101100100100000011100001001011001011110001010011010101111001;  // -1960571374 -876268167
      11'h513: T=64'b1000101100111000100110011100011011001011100101110101010110001010;  // -1959224890 -879274614
      11'h514: T=64'b1000101101001101001101110111110111001011011010010111110110110001;  // -1957873795 -882278991
      11'h515: T=64'b1000101101100001111001110011001111001011001110111010110111110011;  // -1956518093 -885281293
      11'h516: T=64'b1000101101110110101010001110010111001011000011011110011001011001;  // -1955157787 -888281511
      11'h517: T=64'b1000101110001011011111001001000011001010111000000010011011101000;  // -1953792880 -891279640
      11'h518: T=64'b1000101110100000011000100011000011001010101100100110111110101010;  // -1952423376 -894275670
      11'h519: T=64'b1000101110110101010110011100001011001010100001001100000010100011;  // -1951049278 -897269597
      11'h51a: T=64'b1000101111001010011000110100010011001010010101110001100111011100;  // -1949670588 -900261412
      11'h51b: T=64'b1000101111011111011111101011000111001010001010010111101101011011;  // -1948287311 -903251109
      11'h51c: T=64'b1000101111110100101011000000011011001001111110111110010100100111;  // -1946899450 -906238681
      11'h51d: T=64'b1000110000001001111010110100000111001001110011100101011101001000;  // -1945507007 -909224120
      11'h51e: T=64'b1000110000011111001111000101111011001001101000001101000111000101;  // -1944109986 -912207419
      11'h51f: T=64'b1000110000110100100111110101100111001001011100110101010010100100;  // -1942708391 -915188572
      11'h520: T=64'b1000110001001010000101000011000011001001010001011101111111101101;  // -1941302224 -918167571
      11'h521: T=64'b1000110001011111100110101101111111001001000110000111001110100110;  // -1939891489 -921144410
      11'h522: T=64'b1000110001110101001100110110001111001000111010110000111111010110;  // -1938476189 -924119082
      11'h523: T=64'b1000110010001010110111011011100011001000101111011011010010000110;  // -1937056328 -927091578
      11'h524: T=64'b1000110010100000100110011101101111001000100100000110000110111010;  // -1935631909 -930061894
      11'h525: T=64'b1000110010110110011001111100100111001000011000110001011101111100;  // -1934202935 -933030020
      11'h526: T=64'b1000110011001100010001110111111011001000001101011101010111010000;  // -1932769410 -935995952
      11'h527: T=64'b1000110011100010001110001111011111001000000010001001110011000000;  // -1931331337 -938959680
      11'h528: T=64'b1000110011111000001111000011000111000111110110110110110001010000;  // -1929888719 -941921200
      11'h529: T=64'b1000110100001110010100010010100011000111101011100100010010001010;  // -1928441560 -944880502
      11'h52a: T=64'b1000110100100100011101111101100111000111100000010010010101110010;  // -1926989863 -947837582
      11'h52b: T=64'b1000110100111010101100000100000011000111010101000000111100010001;  // -1925533632 -950792431
      11'h52c: T=64'b1000110101010000111110100101101011000111001001110000000101101101;  // -1924072870 -953745043
      11'h52d: T=64'b1000110101100111010101100010010011000110111110011111110010001110;  // -1922607580 -956695410
      11'h52e: T=64'b1000110101111101110000111001101011000110110011010000000001111001;  // -1921137766 -959643527
      11'h52f: T=64'b1000110110010100010000101011100011000110101000000000110100110111;  // -1919663432 -962589385
      11'h530: T=64'b1000110110101010110100110111110011000110011100110010001011001110;  // -1918184580 -965532978
      11'h531: T=64'b1000110111000001011101011110000111000110010001100100000101000101;  // -1916701215 -968474299
      11'h532: T=64'b1000110111011000001010011110010111000110000110010110100010100011;  // -1915213339 -971413341
      11'h533: T=64'b1000110111101110111011111000001111000101111011001001100011101110;  // -1913720957 -974350098
      11'h534: T=64'b1000111000000101110001101011100011000101101111111101001000101111;  // -1912224072 -977284561
      11'h535: T=64'b1000111000011100101011111000000111000101100100110001010001101011;  // -1910722687 -980216725
      11'h536: T=64'b1000111000110011101010011101101011000101011001100101111110101001;  // -1909216806 -983146583
      11'h537: T=64'b1000111001001010101101011100000011000101001110011011001111110001;  // -1907706432 -986074127
      11'h538: T=64'b1000111001100001110100110010111111000101000011010001000101001001;  // -1906191569 -988999351
      11'h539: T=64'b1000111001111001000000100010001111000100111000000111011110111001;  // -1904672221 -991922247
      11'h53a: T=64'b1000111010010000010000101001100111000100101100111110011101000111;  // -1903148391 -994842809
      11'h53b: T=64'b1000111010100111100101001000110111000100100001110101111111111001;  // -1901620083 -997761031
      11'h53c: T=64'b1000111010111110111101111111110011000100010110101110000111010111;  // -1900087300 -1000676905
      11'h53d: T=64'b1000111011010110011011001110001011000100001011100110110011101001;  // -1898550046 -1003590423
      11'h53e: T=64'b1000111011101101111100110011110011000100000000100000000100110011;  // -1897008324 -1006501581
      11'h53f: T=64'b1000111100000101100010110000010111000011110101011001111010111110;  // -1895462139 -1009410370
      11'h540: T=64'b1000111100011101001101000011101111000011101010010100010110010000;  // -1893911493 -1012316784
      11'h541: T=64'b1000111100110100111011101101100111000011011111001111010110110001;  // -1892356391 -1015220815
      11'h542: T=64'b1000111101001100101110101101110011000011010100001010111100100110;  // -1890796836 -1018122458
      11'h543: T=64'b1000111101100100100110000100000011000011001001000111000111110111;  // -1889232832 -1021021705
      11'h544: T=64'b1000111101111100100001110000001011000010111110000011111000101011;  // -1887664382 -1023918549
      11'h545: T=64'b1000111110010100100001110001111011000010110011000001001111000111;  // -1886091490 -1026812985
      11'h546: T=64'b1000111110101100100110001001000011000010100111111111001011010101;  // -1884514160 -1029705003
      11'h547: T=64'b1000111111000100101110110101010011000010011100111101101101011001;  // -1882932396 -1032594599
      11'h548: T=64'b1000111111011100111011110110011111000010010001111100110101011011;  // -1881346201 -1035481765
      11'h549: T=64'b1000111111110101001101001100010111000010000110111100100011100001;  // -1879755579 -1038366495
      11'h54a: T=64'b1001000000001101100010110110101011000001111011111100110111110011;  // -1878160534 -1041248781
      11'h54b: T=64'b1001000000100101111100110101001111000001110000111101110010010111;  // -1876561069 -1044128617
      11'h54c: T=64'b1001000000111110011011000111110011000001100101111111010011010100;  // -1874957188 -1047005996
      11'h54d: T=64'b1001000001010110111101101110000011000001011011000001011010110001;  // -1873348896 -1049880911
      11'h54e: T=64'b1001000001101111100100100111110111000001010000000100001000110100;  // -1871736195 -1052753356
      11'h54f: T=64'b1001000010001000001111110100111011000001000101000111011101100100;  // -1870119090 -1055623324
      11'h550: T=64'b1001000010100000111111010100111111000000111010001011011001001001;  // -1868497585 -1058490807
      11'h551: T=64'b1001000010111001110011000111110111000000101111001111111011101000;  // -1866871683 -1061355800
      11'h552: T=64'b1001000011010010101011001101010111000000100100010101000101001000;  // -1865241387 -1064218296
      11'h553: T=64'b1001000011101011100111100101000111000000011001011010110101110001;  // -1863606703 -1067078287
      11'h554: T=64'b1001000100000100101000001110111111000000001110100001001101101001;  // -1861967633 -1069935767
      11'h555: T=64'b1001000100011101101101001010101011000000000011101000001100110110;  // -1860324182 -1072790730
      11'h556: T=64'b1001000100110110110110010111111010111111111000101111110011100000;  // -1858676354 -1075643168
      11'h557: T=64'b1001000101010000000011110110100010111111101101111000000001101101;  // -1857024152 -1078493075
      11'h558: T=64'b1001000101101001010101100110010010111111100011000000110111100011;  // -1855367580 -1081340445
      11'h559: T=64'b1001000110000010101011100110111010111111011000001010010101001010;  // -1853706642 -1084185270
      11'h55a: T=64'b1001000110011100000101111000000110111111001101010100011010101001;  // -1852041343 -1087027543
      11'h55b: T=64'b1001000110110101100100011001101110111111000010011111001000000101;  // -1850371685 -1089867259
      11'h55c: T=64'b1001000111001111000111001011011110111110110111101010011101100110;  // -1848697673 -1092704410
      11'h55d: T=64'b1001000111101000101110001101000110111110101100110110011011010010;  // -1847019311 -1095538990
      11'h55e: T=64'b1001001000000010011001011110010110111110100010000011000001010000;  // -1845336603 -1098370992
      11'h55f: T=64'b1001001000011100001000111111000010111110010111010000001111100110;  // -1843649552 -1101200410
      11'h560: T=64'b1001001000110101111100101110110010111110001100011110000110011100;  // -1841958164 -1104027236
      11'h561: T=64'b1001001001001111110100101101100010111110000001101100100101111000;  // -1840262440 -1106851464
      11'h562: T=64'b1001001001101001110000111010110110111101110110111011101110000000;  // -1838562387 -1109673088
      11'h563: T=64'b1001001010000011110001010110100110111101101100001011011110111011;  // -1836858007 -1112492101
      11'h564: T=64'b1001001010011101110110000000011110111101100001011011111000110000;  // -1835149305 -1115308496
      11'h565: T=64'b1001001010110111111110111000001110111101010110101100111011100110;  // -1833436285 -1118122266
      11'h566: T=64'b1001001011010010001011111101100110111101001011111110100111100010;  // -1831718951 -1120933406
      11'h567: T=64'b1001001011101100011101010000011010111101000001010000111100101101;  // -1829997306 -1123741907
      11'h568: T=64'b1001001100000110110010110000010110111100110110100011111011001011;  // -1828271355 -1126547765
      11'h569: T=64'b1001001100100001001100011101001010111100101011110111100011000100;  // -1826541102 -1129350972
      11'h56a: T=64'b1001001100111011101010010110100110111100100001001011110100011111;  // -1824806551 -1132151521
      11'h56b: T=64'b1001001101010110001100011100011010111100010110100000101111100010;  // -1823067706 -1134949406
      11'h56c: T=64'b1001001101110000110010101110010110111100001011110110010100010100;  // -1821324571 -1137744620
      11'h56d: T=64'b1001001110001011011101001100000110111100000001001100100010111011;  // -1819577151 -1140537157
      11'h56e: T=64'b1001001110100110001011110101100010111011110110100011011011011101;  // -1817825448 -1143327011
      11'h56f: T=64'b1001001111000000111110101010001110111011101011111010111110000010;  // -1816069469 -1146114174
      11'h570: T=64'b1001001111011011110101101010000110111011100001010011001010110000;  // -1814309215 -1148898640
      11'h571: T=64'b1001001111110110110000110100101110111011010110101100000001101101;  // -1812544693 -1151680403
      11'h572: T=64'b1001010000010001110000001001111010111011001100000101100011000001;  // -1810775906 -1154459455
      11'h573: T=64'b1001010000101100110011101001011110111011000001011111101110110001;  // -1809002857 -1157235791
      11'h574: T=64'b1001010001000111111011010011000010111010110110111010100101000100;  // -1807225552 -1160009404
      11'h575: T=64'b1001010001100011000111000110011010111010101100010110000110000000;  // -1805443994 -1162780288
      11'h576: T=64'b1001010001111110010111000011010010111010100001110010010001101101;  // -1803658188 -1165548435
      11'h577: T=64'b1001010010011001101011001001011010111010010111001111001000010001;  // -1801868138 -1168313839
      11'h578: T=64'b1001010010110101000011011000100010111010001100101100101001110001;  // -1800073848 -1171076495
      11'h579: T=64'b1001010011010000011111110000011010111010000010001010110110010101;  // -1798275322 -1173836395
      11'h57a: T=64'b1001010011101100000000010000110010111001110111101001101110000100;  // -1796472564 -1176593532
      11'h57b: T=64'b1001010100000111100100111001010110111001101101001001010001000011;  // -1794665579 -1179347901
      11'h57c: T=64'b1001010100100011001101101001110010111001100010101001011111011001;  // -1792854372 -1182099495
      11'h57d: T=64'b1001010100111110111010100001111110111001011000001010011001001100;  // -1791038945 -1184848308
      11'h57e: T=64'b1001010101011010101011100001100010111001001101101011111110100100;  // -1789219304 -1187594332
      11'h57f: T=64'b1001010101110110100000101000001110111001000011001110001111100111;  // -1787395453 -1190337561
      11'h580: T=64'b1001010110010010011001110101110110111000111000110001001100011010;  // -1785567395 -1193077990
      11'h581: T=64'b1001010110101110010111001001111110111000101110010100110101000101;  // -1783735137 -1195815611
      11'h582: T=64'b1001010111001010011000100100100010111000100011111001001001101101;  // -1781898680 -1198550419
      11'h583: T=64'b1001010111100110011110000101000110111000011001011110001010011010;  // -1780058031 -1201282406
      11'h584: T=64'b1001011000000010100111101011011010111000001111000011110111010010;  // -1778213194 -1204011566
      11'h585: T=64'b1001011000011110110101010111010010111000000100101010010000011010;  // -1776364172 -1206737894
      11'h586: T=64'b1001011000111011000111001000011010110111111010010001010101111011;  // -1774510970 -1209461381
      11'h587: T=64'b1001011001010111011100111110100010110111101111111001000111111001;  // -1772653592 -1212182023
      11'h588: T=64'b1001011001110011110110111001010110110111100101100001100110011100;  // -1770792043 -1214899812
      11'h589: T=64'b1001011010010000010100111000100010110111011011001010110001101001;  // -1768926328 -1217614743
      11'h58a: T=64'b1001011010101100110110111011111110110111010000110100101001101000;  // -1767056449 -1220326808
      11'h58b: T=64'b1001011011001001011101000011001110110111000110011111001110011110;  // -1765182413 -1223036002
      11'h58c: T=64'b1001011011100110000111001110000110110110111100001010100000010010;  // -1763304223 -1225742318
      11'h58d: T=64'b1001011100000010110101011100010010110110110001110110011111001011;  // -1761421884 -1228445749
      11'h58e: T=64'b1001011100011111100111101101011110110110100111100011001011001110;  // -1759535401 -1231146290
      11'h58f: T=64'b1001011100111100011110000001100010110110011101010000100100100010;  // -1757644776 -1233843934
      11'h590: T=64'b1001011101011001011000011000000010110110010010111110101011001101;  // -1755750016 -1236538675
      11'h591: T=64'b1001011101110110010110110000101110110110001000101101011111010110;  // -1753851125 -1239230506
      11'h592: T=64'b1001011110010011011001001011011010110101111110011101000001000011;  // -1751948106 -1241919421
      11'h593: T=64'b1001011110110000011111100111101110110101110100001101010000011011;  // -1750040965 -1244605413
      11'h594: T=64'b1001011111001101101010000101011010110101101001111110001101100011;  // -1748129706 -1247288477
      11'h595: T=64'b1001011111101010111000100100001010110101011111101111111000100010;  // -1746214334 -1249968606
      11'h596: T=64'b1001100000001000001011000011110010110101010101100010010001011111;  // -1744294852 -1252645793
      11'h597: T=64'b1001100000100101100001100011111010110101001011010101011000011111;  // -1742371266 -1255320033
      11'h598: T=64'b1001100001000010111100000100010010110101000001001001001101101001;  // -1740443580 -1257991319
      11'h599: T=64'b1001100001100000011010100100101010110100110110111101110001000011;  // -1738511798 -1260659645
      11'h59a: T=64'b1001100001111101111101000100101010110100101100110011000010110011;  // -1736575926 -1263325005
      11'h59b: T=64'b1001100010011011100011100100000110110100100010101001000011000001;  // -1734635967 -1265987391
      11'h59c: T=64'b1001100010111001001110000010100110110100011000011111110001110001;  // -1732691927 -1268646799
      11'h59d: T=64'b1001100011010110111100011111111110110100001110010111001111001010;  // -1730743809 -1271303222
      11'h59e: T=64'b1001100011110100101110111011110110110100000100001111011011010100;  // -1728791619 -1273956652
      11'h59f: T=64'b1001100100010010100101010101111110110011111010001000010110010010;  // -1726835361 -1276607086
      11'h5a0: T=64'b1001100100110000011111101110000110110011110000000010000000001101;  // -1724875039 -1279254515
      11'h5a1: T=64'b1001100101001110011110000011110110110011100101111100011001001010;  // -1722910659 -1281898934
      11'h5a2: T=64'b1001100101101100100000010111000010110011011011110111100001001111;  // -1720942224 -1284540337
      11'h5a3: T=64'b1001100110001010100110100111010010110011010001110011011000100011;  // -1718969740 -1287178717
      11'h5a4: T=64'b1001100110101000110000110100010110110011000111101111111111001100;  // -1716993211 -1289814068
      11'h5a5: T=64'b1001100111000110111110111101111110110010111101101101010101010000;  // -1715012641 -1292446384
      11'h5a6: T=64'b1001100111100101010001000011110010110010110011101011011010110110;  // -1713028036 -1295075658
      11'h5a7: T=64'b1001101000000011100111000101100010110010101001101010010000000010;  // -1711039400 -1297701886
      11'h5a8: T=64'b1001101000100010000001000010111010110010011111101001110100111101;  // -1709046738 -1300325059
      11'h5a9: T=64'b1001101001000000011110111011100110110010010101101010001001101011;  // -1707050055 -1302945173
      11'h5aa: T=64'b1001101001011111000000101111011010110010001011101011001110010011;  // -1705049354 -1305562221
      11'h5ab: T=64'b1001101001111101100110011101111010110010000001101101000010111011;  // -1703044642 -1308176197
      11'h5ac: T=64'b1001101010011100010000000110111110110001110111101111100111101001;  // -1701035921 -1310787095
      11'h5ad: T=64'b1001101010111010111101101010000110110001101101110010111100100100;  // -1699023199 -1313394908
      11'h5ae: T=64'b1001101011011001101111000111001010110001100011110111000001110001;  // -1697006478 -1315999631
      11'h5af: T=64'b1001101011111000100100011101110010110001011001111011110111010111;  // -1694985764 -1318601257
      11'h5b0: T=64'b1001101100010111011101101101101110110001010000000001011101011100;  // -1692961061 -1321199780
      11'h5b1: T=64'b1001101100110110011010110110100110110001000110000111110100000110;  // -1690932375 -1323795194
      11'h5b2: T=64'b1001101101010101011011111000001010110000111100001110111011011011;  // -1688899710 -1326387493
      11'h5b3: T=64'b1001101101110100100000110010000110110000110010010110110011100000;  // -1686863071 -1328976672
      11'h5b4: T=64'b1001101110010011101001100100000110110000101000011111011100011110;  // -1684822463 -1331562722
      11'h5b5: T=64'b1001101110110010110110001101111110110000011110101000110110011000;  // -1682777889 -1334145640
      11'h5b6: T=64'b1001101111010010000110101111001110110000010100110011000001010110;  // -1680729357 -1336725418
      11'h5b7: T=64'b1001101111110001011011000111101110110000001010111101111101011101;  // -1678676869 -1339302051
      11'h5b8: T=64'b1001110000010000110011010111000110110000000001001001101010110100;  // -1676620431 -1341875532
      11'h5b9: T=64'b1001110000110000001111011101000010101111110111010110001001100000;  // -1674560048 -1344445856
      11'h5ba: T=64'b1001110001001111101111011001010010101111101101100011011001101000;  // -1672495724 -1347013016
      11'h5bb: T=64'b1001110001101111010011001011011110101111100011110001011011010001;  // -1670427465 -1349577007
      11'h5bc: T=64'b1001110010001110111010110011010010101111011010000000001110100010;  // -1668355276 -1352137822
      11'h5bd: T=64'b1001110010101110100110010000100010101111010000001111110011100001;  // -1666279160 -1354695455
      11'h5be: T=64'b1001110011001110010101100010110010101111000110100000001010010100;  // -1664199124 -1357249900
      11'h5bf: T=64'b1001110011101110001000101001110110101110111100110001010011000000;  // -1662115171 -1359801152
      11'h5c0: T=64'b1001110100001101111111100101010010101110110011000011001101101100;  // -1660027308 -1362349204
      11'h5c1: T=64'b1001110100101101111010010100111010101110101001010101111010011110;  // -1657935538 -1364894050
      11'h5c2: T=64'b1001110101001101111000111000010110101110011111101001011001011100;  // -1655839867 -1367435684
      11'h5c3: T=64'b1001110101101101111011001111010110101110010101111101101010101011;  // -1653740299 -1369974101
      11'h5c4: T=64'b1001110110001110000001011001100010101110001100010010101110010010;  // -1651636840 -1372509294
      11'h5c5: T=64'b1001110110101110001011010110100110101110000010101000100100010111;  // -1649529495 -1375041257
      11'h5c6: T=64'b1001110111001110011001000110010010101101111000111111001100111111;  // -1647418268 -1377569985
      11'h5c7: T=64'b1001110111101110101010101000001110101101101111010110101000010001;  // -1645303165 -1380095471
      11'h5c8: T=64'b1001111000001110111111111100001010101101100101101110110110010010;  // -1643184190 -1382617710
      11'h5c9: T=64'b1001111000101111011001000001101110101101011100000111110111001001;  // -1641061349 -1385136695
      11'h5ca: T=64'b1001111001001111110101111000101010101101010010100001101010111011;  // -1638934646 -1387652421
      11'h5cb: T=64'b1001111001110000010110100000101010101101001000111100010001101110;  // -1636804086 -1390164882
      11'h5cc: T=64'b1001111010010000111010111001010110101100111111010111101011101001;  // -1634669675 -1392674071
      11'h5cd: T=64'b1001111010110001100011000010011110101100110101110011111000110001;  // -1632531417 -1395179983
      11'h5ce: T=64'b1001111011010010001110111011101010101100101100010000111001001011;  // -1630389318 -1397682613
      11'h5cf: T=64'b1001111011110010111110100100101010101100100010101110101100111111;  // -1628243382 -1400181953
      11'h5d0: T=64'b1001111100010011110001111101000110101100011001001101010100010001;  // -1626093615 -1402677999
      11'h5d1: T=64'b1001111100110100101001000100101010101100001111101100101111001000;  // -1623940022 -1405170744
      11'h5d2: T=64'b1001111101010101100011111011000110101100000110001100111101101001;  // -1621782607 -1407660183
      11'h5d3: T=64'b1001111101110110100010100000000010101011111100101101111111111011;  // -1619621376 -1410146309
      11'h5d4: T=64'b1001111110010111100100110011001010101011110011001111110110000011;  // -1617456334 -1412629117
      11'h5d5: T=64'b1001111110111000101010110100001010101011101001110010100000000111;  // -1615287486 -1415108601
      11'h5d6: T=64'b1001111111011001110100100010101110101011100000010101111110001101;  // -1613114837 -1417584755
      11'h5d7: T=64'b1001111111111011000001111110100010101011010110111010010000011011;  // -1610938392 -1420057573
      11'h5d8: T=64'b1010000000011100010011000111001110101011001101011111010110110110;  // -1608758157 -1422527050
      11'h5d9: T=64'b1010000000111101100111111100100010101011000100000101010001100101;  // -1606574136 -1424993179
      11'h5da: T=64'b1010000001011111000000011110001010101010111010101100000000101100;  // -1604386334 -1427455956
      11'h5db: T=64'b1010000010000000011100101011101110101010110001010011100100010011;  // -1602194757 -1429915373
      11'h5dc: T=64'b1010000010100001111100100100111010101010100111111011111100011110;  // -1599999410 -1432371426
      11'h5dd: T=64'b1010000011000011100000001001011010101010011110100101001001010100;  // -1597800298 -1434824108
      11'h5de: T=64'b1010000011100101000111011000110110101010010101001111001010111010;  // -1595597427 -1437273414
      11'h5df: T=64'b1010000100000110110010010010111110101010001011111010000001010110;  // -1593390801 -1439719338
      11'h5e0: T=64'b1010000100101000100000110111011110101010000010100101101100101110;  // -1591180425 -1442161874
      11'h5e1: T=64'b1010000101001010010011000101111110101001111001010010001101001000;  // -1588966305 -1444601016
      11'h5e2: T=64'b1010000101101100001000111110001010101001101111111111100010101001;  // -1586748446 -1447036759
      11'h5e3: T=64'b1010000110001110000010011111101010101001100110101101101101010111;  // -1584526854 -1449469097
      11'h5e4: T=64'b1010000110101111111111101010001110101001011101011100101101010111;  // -1582301533 -1451898025
      11'h5e5: T=64'b1010000111010010000000011101100010101001010100001100100010110000;  // -1580072488 -1454323536
      11'h5e6: T=64'b1010000111110100000100111001001010101001001010111101001101100111;  // -1577839726 -1456745625
      11'h5e7: T=64'b1010001000010110001100111100111010101001000001101110101110000010;  // -1575603250 -1459164286
      11'h5e8: T=64'b1010001000111000011000101000010110101000111000100001000100000111;  // -1573363067 -1461579513
      11'h5e9: T=64'b1010001001011010100111111011001010101000101111010100001111111011;  // -1571119182 -1463991301
      11'h5ea: T=64'b1010001001111100111010110101000010101000100110001000010001100100;  // -1568871600 -1466399644
      11'h5eb: T=64'b1010001010011111010001010101101010101000011100111101001001000111;  // -1566620326 -1468804537
      11'h5ec: T=64'b1010001011000001101011011100101010101000010011110010110110101011;  // -1564365366 -1471205973
      11'h5ed: T=64'b1010001011100100001001001001101110101000001010101001011010010100;  // -1562106725 -1473603948
      11'h5ee: T=64'b1010001100000110101010011100100110101000000001100000110100001001;  // -1559844407 -1475998455
      11'h5ef: T=64'b1010001100101001001111010100110010100111111000011001000100001111;  // -1557578420 -1478389489
      11'h5f0: T=64'b1010001101001011110111110010000110100111101111010010001010101100;  // -1555308767 -1480777044
      11'h5f1: T=64'b1010001101101110100011110100001010100111100110001100000111100110;  // -1553035454 -1483161114
      11'h5f2: T=64'b1010001110010001010011011010100010100111011101000110111011000001;  // -1550758488 -1485541695
      11'h5f3: T=64'b1010001110110100000110100101000110100111010100000010100101000100;  // -1548477871 -1487918780
      11'h5f4: T=64'b1010001111010110111101010011010010100111001010111111000101110100;  // -1546193612 -1490292364
      11'h5f5: T=64'b1010001111111001110111100100111010100111000001111100011101010111;  // -1543905714 -1492662441
      11'h5f6: T=64'b1010010000011100110101011001101010100110111000111010101011110011;  // -1541614182 -1495029005
      11'h5f7: T=64'b1010010000111111110110110001000010100110101111111001110001001100;  // -1539319024 -1497392052
      11'h5f8: T=64'b1010010001100010111011101010110110100110100110111001101101101001;  // -1537020243 -1499751575
      11'h5f9: T=64'b1010010010000110000100000110101110100110011101111010100001001111;  // -1534717845 -1502107569
      11'h5fa: T=64'b1010010010101001010000000100010010100110010100111100001100000011;  // -1532411836 -1504460029
      11'h5fb: T=64'b1010010011001100011111100011001010100110001011111110101110001100;  // -1530102222 -1506808948
      11'h5fc: T=64'b1010010011101111110010100011001010100110000011000010000111101110;  // -1527789006 -1509154322
      11'h5fd: T=64'b1010010100010011001001000011110010100101111010000110011000110000;  // -1525472196 -1511496144
      11'h5fe: T=64'b1010010100110110100011000100110010100101110001001011100001010110;  // -1523151796 -1513834410
      11'h5ff: T=64'b1010010101011010000000100101110010100101101000010001100001100111;  // -1520827812 -1516169113
      11'h600: T=64'b1010010101111101100001100110011110100101011111011000011001100111;  // -1518500249 -1518500249
      11'h601: T=64'b1010010110100001000110000110011110100101010110100000001001011100;  // -1516169113 -1520827812
      11'h602: T=64'b1010010111000100101110000101011010100101001101101000110001001100;  // -1513834410 -1523151796
      11'h603: T=64'b1010010111101000011001100011000010100101000100110010010000111100;  // -1511496144 -1525472196
      11'h604: T=64'b1010011000001100001000011110111010100100111011111100101000110010;  // -1509154322 -1527789006
      11'h605: T=64'b1010011000101111111010111000110010100100110011000111111000110010;  // -1506808948 -1530102222
      11'h606: T=64'b1010011001010011110000110000001110100100101010010100000001000100;  // -1504460029 -1532411836
      11'h607: T=64'b1010011001110111101010000100111110100100100001100001000001101011;  // -1502107569 -1534717845
      11'h608: T=64'b1010011010011011100110110110100110100100011000101110111010101101;  // -1499751575 -1537020243
      11'h609: T=64'b1010011010111111100111000100110010100100001111111101101100010000;  // -1497392052 -1539319024
      11'h60a: T=64'b1010011011100011101010101111001110100100000111001101010110011010;  // -1495029005 -1541614182
      11'h60b: T=64'b1010011100000111110001110101011110100011111110011101111001001110;  // -1492662441 -1543905714
      11'h60c: T=64'b1010011100101011111100010111010010100011110101101111010100110100;  // -1490292364 -1546193612
      11'h60d: T=64'b1010011101010000001010010100010010100011101101000001101001010001;  // -1487918780 -1548477871
      11'h60e: T=64'b1010011101110100011011101100000110100011100100010100110110101000;  // -1485541695 -1550758488
      11'h60f: T=64'b1010011110011000110000011110011010100011011011101000111101000010;  // -1483161114 -1553035454
      11'h610: T=64'b1010011110111101001000101010110010100011010010111101111100100001;  // -1480777044 -1555308767
      11'h611: T=64'b1010011111100001100100010000111110100011001010010011110101001100;  // -1478389489 -1557578420
      11'h612: T=64'b1010100000000110000011010000100110100011000001101010100111001001;  // -1475998455 -1559844407
      11'h613: T=64'b1010100000101010100101101001010010100010111001000010010010011011;  // -1473603948 -1562106725
      11'h614: T=64'b1010100001001111001011011010101110100010110000011010110111001010;  // -1471205973 -1564365366
      11'h615: T=64'b1010100001110011110100100100011110100010100111110100010101011010;  // -1468804537 -1566620326
      11'h616: T=64'b1010100010011000100001000110010010100010011111001110101101010000;  // -1466399644 -1568871600
      11'h617: T=64'b1010100010111101010000111111101110100010010110101001111110110010;  // -1463991301 -1571119182
      11'h618: T=64'b1010100011100010000100010000011110100010001110000110001010000101;  // -1461579513 -1573363067
      11'h619: T=64'b1010100100000110111010111000001010100010000101100011001111001110;  // -1459164286 -1575603250
      11'h61a: T=64'b1010100100101011110100110110011110100001111101000001001110010010;  // -1456745625 -1577839726
      11'h61b: T=64'b1010100101010000110010001011000010100001110100100000000111011000;  // -1454323536 -1580072488
      11'h61c: T=64'b1010100101110101110010110101011110100001101011111111111010100011;  // -1451898025 -1582301533
      11'h61d: T=64'b1010100110011010110110110101011110100001100011100000100111111010;  // -1449469097 -1584526854
      11'h61e: T=64'b1010100110111111111110001010100110100001011011000010001111100010;  // -1447036759 -1586748446
      11'h61f: T=64'b1010100111100101001000110100100010100001010010100100110001011111;  // -1444601016 -1588966305
      11'h620: T=64'b1010101000001010010110110010111010100001001010001000001101110111;  // -1442161874 -1591180425
      11'h621: T=64'b1010101000101111101000000101011010100001000001101100100100101111;  // -1439719338 -1593390801
      11'h622: T=64'b1010101001010100111100101011101010100000111001010001110110001101;  // -1437273414 -1595597427
      11'h623: T=64'b1010101001111010010100100101010010100000110000111000000010010110;  // -1434824108 -1597800298
      11'h624: T=64'b1010101010011111101111110001111010100000101000011111001001001110;  // -1432371426 -1599999410
      11'h625: T=64'b1010101011000101001110010001001110100000100000000111001010111011;  // -1429915373 -1602194757
      11'h626: T=64'b1010101011101010110000000010110010100000010111110000000111100010;  // -1427455956 -1604386334
      11'h627: T=64'b1010101100010000010101000110010110100000001111011001111111001000;  // -1424993179 -1606574136
      11'h628: T=64'b1010101100110101111101011011011010100000000111000100110001110011;  // -1422527050 -1608758157
      11'h629: T=64'b1010101101011011101001000001101110011111111110110000011111101000;  // -1420057573 -1610938392
      11'h62a: T=64'b1010101110000001010111111000110110011111110110011101001000101011;  // -1417584755 -1613114837
      11'h62b: T=64'b1010101110100111001010000000011110011111101110001010101101000010;  // -1415108601 -1615287486
      11'h62c: T=64'b1010101111001100111111011000001110011111100101111001001100110010;  // -1412629117 -1617456334
      11'h62d: T=64'b1010101111110010110111111111101110011111011101101000101000000000;  // -1410146309 -1619621376
      11'h62e: T=64'b1010110000011000110011110110100110011111010101011000111110110001;  // -1407660183 -1621782607
      11'h62f: T=64'b1010110000111110110010111100100010011111001101001010010001001010;  // -1405170744 -1623940022
      11'h630: T=64'b1010110001100100110101010001000110011111000100111100011111010001;  // -1402677999 -1626093615
      11'h631: T=64'b1010110010001010111010110011111110011110111100101111101001001010;  // -1400181953 -1628243382
      11'h632: T=64'b1010110010110001000011100100101110011110110100100011101110111010;  // -1397682613 -1630389318
      11'h633: T=64'b1010110011010111001111100011000110011110101100011000110000100111;  // -1395179983 -1632531417
      11'h634: T=64'b1010110011111101011110101110100110011110100100001110101110010101;  // -1392674071 -1634669675
      11'h635: T=64'b1010110100100011110001000110111010011110011100000101101000001010;  // -1390164882 -1636804086
      11'h636: T=64'b1010110101001010000110101011101110011110010011111101011110001010;  // -1387652421 -1638934646
      11'h637: T=64'b1010110101110000011111011100100110011110001011110110010000011011;  // -1385136695 -1641061349
      11'h638: T=64'b1010110110010110111011011001001010011110000011101111111111000010;  // -1382617710 -1643184190
      11'h639: T=64'b1010110110111101011010100001000110011101111011101010101010000011;  // -1380095471 -1645303165
      11'h63a: T=64'b1010110111100011111100110011111110011101110011100110010001100100;  // -1377569985 -1647418268
      11'h63b: T=64'b1010111000001010100010010001011110011101101011100010110101101001;  // -1375041257 -1649529495
      11'h63c: T=64'b1010111000110001001010111001001010011101100011100000010110011000;  // -1372509294 -1651636840
      11'h63d: T=64'b1010111001010111110110101010101110011101011011011110110011110101;  // -1369974101 -1653740299
      11'h63e: T=64'b1010111001111110100101100101110010011101010011011110001110000101;  // -1367435684 -1655839867
      11'h63f: T=64'b1010111010100101010111101001111010011101001011011110100101001110;  // -1364894050 -1657935538
      11'h640: T=64'b1010111011001100001100110110110010011101000011011111111001010100;  // -1362349204 -1660027308
      11'h641: T=64'b1010111011110011000101001100000010011100111011100010001010011101;  // -1359801152 -1662115171
      11'h642: T=64'b1010111100011010000000101001010010011100110011100101011000101100;  // -1357249900 -1664199124
      11'h643: T=64'b1010111101000000111111001110000110011100101011101001100100001000;  // -1354695455 -1666279160
      11'h644: T=64'b1010111101101000000000111010001010011100100011101110101100110100;  // -1352137822 -1668355276
      11'h645: T=64'b1010111110001111000101101101000110011100011011110100110010110111;  // -1349577007 -1670427465
      11'h646: T=64'b1010111110110110001101100110100010011100010011111011110110010100;  // -1347013016 -1672495724
      11'h647: T=64'b1010111111011101011000100110000010011100001100000011110111010000;  // -1344445856 -1674560048
      11'h648: T=64'b1011000000000100100110101011010010011100000100001100110101110001;  // -1341875532 -1676620431
      11'h649: T=64'b1011000000101011110111110101110110011011111100010110110001111011;  // -1339302051 -1678676869
      11'h64a: T=64'b1011000001010011001100000101011010011011110100100001101011110011;  // -1336725418 -1680729357
      11'h64b: T=64'b1011000001111010100011011001100010011011101100101101100011011111;  // -1334145640 -1682777889
      11'h64c: T=64'b1011000010100001111101110001111010011011100100111010011001000001;  // -1331562722 -1684822463
      11'h64d: T=64'b1011000011001001011011001110000010011011011101001000001100100001;  // -1328976672 -1686863071
      11'h64e: T=64'b1011000011110000111011101101101110011011010101010110111110000010;  // -1326387493 -1688899710
      11'h64f: T=64'b1011000100011000011111010000011010011011001101100110101101101001;  // -1323795194 -1690932375
      11'h650: T=64'b1011000101000000000101110101110010011011000101110111011011011011;  // -1321199780 -1692961061
      11'h651: T=64'b1011000101100111101111011101011110011010111110001001000111011100;  // -1318601257 -1694985764
      11'h652: T=64'b1011000110001111011100000111000110011010110110011011110001110010;  // -1315999631 -1697006478
      11'h653: T=64'b1011000110110111001011110010010010011010101110101111011010100001;  // -1313394908 -1699023199
      11'h654: T=64'b1011000111011110111110011110100110011010100111000100000001101111;  // -1310787095 -1701035921
      11'h655: T=64'b1011001000000110110100001011101110011010011111011001100111011110;  // -1308176197 -1703044642
      11'h656: T=64'b1011001000101110101100111001001110011010010111110000001011110110;  // -1305562221 -1705049354
      11'h657: T=64'b1011001001010110101000100110101110011010010000000111101110111001;  // -1302945173 -1707050055
      11'h658: T=64'b1011001001111110100111010011110110011010001000100000010000101110;  // -1300325059 -1709046738
      11'h659: T=64'b1011001010100110101001000000001010011010000000111001110001011000;  // -1297701886 -1711039400
      11'h65a: T=64'b1011001011001110101101101011011010011001111001010100010000111100;  // -1295075658 -1713028036
      11'h65b: T=64'b1011001011110110110101010101000010011001110001101111101111011111;  // -1292446384 -1715012641
      11'h65c: T=64'b1011001100011110111111111100110010011001101010001100001101000101;  // -1289814068 -1716993211
      11'h65d: T=64'b1011001101000111001101100010001110011001100010101001101001110100;  // -1287178717 -1718969740
      11'h65e: T=64'b1011001101101111011110000100111110011001011011001000000101110000;  // -1284540337 -1720942224
      11'h65f: T=64'b1011001110010111110001100100101010011001010011100111100000111101;  // -1281898934 -1722910659
      11'h660: T=64'b1011001111000000001000000000110110011001001100000111111011100001;  // -1279254515 -1724875039
      11'h661: T=64'b1011001111101000100001011001001010011001000100101001010101011111;  // -1276607086 -1726835361
      11'h662: T=64'b1011010000010000111101101101010010011000111101001011101110111101;  // -1273956652 -1728791619
      11'h663: T=64'b1011010000111001011100111100101010011000110101101111000111111111;  // -1271303222 -1730743809
      11'h664: T=64'b1011010001100001111111000111000110011000101110010011100000101001;  // -1268646799 -1732691927
      11'h665: T=64'b1011010010001010100100001100000110011000100110111000111001000001;  // -1265987391 -1734635967
      11'h666: T=64'b1011010010110011001100001011001110011000011111011111010001001010;  // -1263325005 -1736575926
      11'h667: T=64'b1011010011011011110111000100001110011000011000000110101001001010;  // -1260659645 -1738511798
      11'h668: T=64'b1011010100000100100100110110100110011000010000101111000001000100;  // -1257991319 -1740443580
      11'h669: T=64'b1011010100101101010101100001111110011000001001011000011000111110;  // -1255320033 -1742371266
      11'h66a: T=64'b1011010101010110001001000101111110011000000010000010110000111100;  // -1252645793 -1744294852
      11'h66b: T=64'b1011010101111110111111100010001010010111111010101110001001000010;  // -1249968606 -1746214334
      11'h66c: T=64'b1011010110100111111000110110001110010111110011011010100001010110;  // -1247288477 -1748129706
      11'h66d: T=64'b1011010111010000110101000001101110010111101100000111111001111011;  // -1244605413 -1750040965
      11'h66e: T=64'b1011010111111001110100000100001110010111100100110110010010110110;  // -1241919421 -1751948106
      11'h66f: T=64'b1011011000100010110101111101011010010111011101100101101100001011;  // -1239230506 -1753851125
      11'h670: T=64'b1011011001001011111010101100110110010111010110010110000110000000;  // -1236538675 -1755750016
      11'h671: T=64'b1011011001110101000010010010001010010111001111000111100000011000;  // -1233843934 -1757644776
      11'h672: T=64'b1011011010011110001100101100111010010111000111111001111011010111;  // -1231146290 -1759535401
      11'h673: T=64'b1011011011000111011001111100101110010111000000101101010111000100;  // -1228445749 -1761421884
      11'h674: T=64'b1011011011110000101010000001001010010110111001100001110011100001;  // -1225742318 -1763304223
      11'h675: T=64'b1011011100011001111100111001111010010110110010010111010000110011;  // -1223036002 -1765182413
      11'h676: T=64'b1011011101000011010010100110100010010110101011001101101110111111;  // -1220326808 -1767056449
      11'h677: T=64'b1011011101101100101011000110100110010110100100000101001110001000;  // -1217614743 -1768926328
      11'h678: T=64'b1011011110010110000110011001110010010110011100111101101110010101;  // -1214899812 -1770792043
      11'h679: T=64'b1011011110111111100100011111100110010110010101110111001111101000;  // -1212182023 -1772653592
      11'h67a: T=64'b1011011111101001000101010111101110010110001110110001110010000110;  // -1209461381 -1774510970
      11'h67b: T=64'b1011100000010010101001000001101010010110000111101101010101110100;  // -1206737894 -1776364172
      11'h67c: T=64'b1011100000111100001111011101001010010110000000101001111010110110;  // -1204011566 -1778213194
      11'h67d: T=64'b1011100001100101111000101001101010010101111001100111100001010001;  // -1201282406 -1780058031
      11'h67e: T=64'b1011100010001111100100100110110110010101110010100110001001001000;  // -1198550419 -1781898680
      11'h67f: T=64'b1011100010111001010011010100010110010101101011100101110010011111;  // -1195815611 -1783735137
      11'h680: T=64'b1011100011100011000100110001101010010101100100100110011101011101;  // -1193077990 -1785567395
      11'h681: T=64'b1011100100001100111000111110011110010101011101101000001010000011;  // -1190337561 -1787395453
      11'h682: T=64'b1011100100110110101111111010010010010101010110101010111000011000;  // -1187594332 -1789219304
      11'h683: T=64'b1011100101100000101001100100110010010101001111101110101000011111;  // -1184848308 -1791038945
      11'h684: T=64'b1011100110001010100101111101100110010101001000110011011010011100;  // -1182099495 -1792854372
      11'h685: T=64'b1011100110110100100101000100001110010101000001111001001110010101;  // -1179347901 -1794665579
      11'h686: T=64'b1011100111011110100110111000010010010100111011000000000100001100;  // -1176593532 -1796472564
      11'h687: T=64'b1011101000001000101011011001010110010100110100000111111100000110;  // -1173836395 -1798275322
      11'h688: T=64'b1011101000110010110010100111000110010100101101010000110110001000;  // -1171076495 -1800073848
      11'h689: T=64'b1011101001011100111100100001000110010100100110011010110010010110;  // -1168313839 -1801868138
      11'h68a: T=64'b1011101010000111001001000110110110010100011111100101110000110100;  // -1165548435 -1803658188
      11'h68b: T=64'b1011101010110001011000011000000010010100011000110001110001100110;  // -1162780288 -1805443994
      11'h68c: T=64'b1011101011011011101010010100010010010100010001111110110100110000;  // -1160009404 -1807225552
      11'h68d: T=64'b1011101100000101111110111011000110010100001011001100111010010111;  // -1157235791 -1809002857
      11'h68e: T=64'b1011101100110000010110001100000110010100000100011100000010011110;  // -1154459455 -1810775906
      11'h68f: T=64'b1011101101011010110000000110110110010011111101101100001101001011;  // -1151680403 -1812544693
      11'h690: T=64'b1011101110000101001100101011000010010011110110111101011010100001;  // -1148898640 -1814309215
      11'h691: T=64'b1011101110101111101011111000001010010011110000001111101010100011;  // -1146114174 -1816069469
      11'h692: T=64'b1011101111011010001101101101110110010011101001100010111101011000;  // -1143327011 -1817825448
      11'h693: T=64'b1011110000000100110010001011101110010011100010110111010011000001;  // -1140537157 -1819577151
      11'h694: T=64'b1011110000101111011001010001010010010011011100001100101011100101;  // -1137744620 -1821324571
      11'h695: T=64'b1011110001011010000010111110001010010011010101100011000111000110;  // -1134949406 -1823067706
      11'h696: T=64'b1011110010000100101111010001111110010011001110111010100101101001;  // -1132151521 -1824806551
      11'h697: T=64'b1011110010101111011110001100010010010011001000010011000111010010;  // -1129350972 -1826541102
      11'h698: T=64'b1011110011011010001111101100101110010011000001101100101100000101;  // -1126547765 -1828271355
      11'h699: T=64'b1011110100000101000011110010110110010010111011000111010100000110;  // -1123741907 -1829997306
      11'h69a: T=64'b1011110100101111111010011110001010010010110100100010111111011001;  // -1120933406 -1831718951
      11'h69b: T=64'b1011110101011010110011101110011010010010101101111111101110000011;  // -1118122266 -1833436285
      11'h69c: T=64'b1011110110000101101111100011000010010010100111011101100000000111;  // -1115308496 -1835149305
      11'h69d: T=64'b1011110110110000101101111011101110010010100000111100010101101001;  // -1112492101 -1836858007
      11'h69e: T=64'b1011110111011011101110111000000010010010011010011100001110101101;  // -1109673088 -1838562387
      11'h69f: T=64'b1011111000000110110010010111100010010010010011111101001011011000;  // -1106851464 -1840262440
      11'h6a0: T=64'b1011111000110001111000011001110010010010001101011111001011101100;  // -1104027236 -1841958164
      11'h6a1: T=64'b1011111001011101000000111110011010010010000111000010001111110000;  // -1101200410 -1843649552
      11'h6a2: T=64'b1011111010001000001100000101000010010010000000100110010111100101;  // -1098370992 -1845336603
      11'h6a3: T=64'b1011111010110011011001101101001010010001111010001011100011010001;  // -1095538990 -1847019311
      11'h6a4: T=64'b1011111011011110101001110110011010010001110011110001110010110111;  // -1092704410 -1848697673
      11'h6a5: T=64'b1011111100001001111100100000010110010001101101011001000110011011;  // -1089867259 -1850371685
      11'h6a6: T=64'b1011111100110101010001101010100110010001100111000001011110000001;  // -1087027543 -1852041343
      11'h6a7: T=64'b1011111101100000101001010100101010010001100000101010111001101110;  // -1084185270 -1853706642
      11'h6a8: T=64'b1011111110001100000011011110001110010001011010010101011001100100;  // -1081340445 -1855367580
      11'h6a9: T=64'b1011111110110111100000000110110110010001010100000000111101101000;  // -1078493075 -1857024152
      11'h6aa: T=64'b1011111111100010111111001110000010010001001101101101100101111110;  // -1075643168 -1858676354
      11'h6ab: T=64'b1100000000001110100000110011011010010001000111011011010010101010;  // -1072790730 -1860324182
      11'h6ac: T=64'b1100000000111010000100110110100110010001000001001010000011101111;  // -1069935767 -1861967633
      11'h6ad: T=64'b1100000001100101101011010111000110010000111010111001111001010001;  // -1067078287 -1863606703
      11'h6ae: T=64'b1100000010010001010100010100100010010000110100101010110011010101;  // -1064218296 -1865241387
      11'h6af: T=64'b1100000010111100111111101110100010010000101110011100110001111101;  // -1061355800 -1866871683
      11'h6b0: T=64'b1100000011101000101101100100100110010000101000001111110101001111;  // -1058490807 -1868497585
      11'h6b1: T=64'b1100000100010100011101110110010010010000100010000011111101001110;  // -1055623324 -1870119090
      11'h6b2: T=64'b1100000101000000010000100011010010010000011011111001001001111101;  // -1052753356 -1871736195
      11'h6b3: T=64'b1100000101101100000101101011000110010000010101101111011011100000;  // -1049880911 -1873348896
      11'h6b4: T=64'b1100000110010111111101001101010010010000001111100110110001111100;  // -1047005996 -1874957188
      11'h6b5: T=64'b1100000111000011110111001001011110010000001001011111001101010011;  // -1044128617 -1876561069
      11'h6b6: T=64'b1100000111101111110011011111001110010000000011011000101101101010;  // -1041248781 -1878160534
      11'h6b7: T=64'b1100001000011011110010001110000110001111111101010011010011000101;  // -1038366495 -1879755579
      11'h6b8: T=64'b1100001001000111110011010101101110001111110111001110111101100111;  // -1035481765 -1881346201
      11'h6b9: T=64'b1100001001110011110110110101100110001111110001001011101101010100;  // -1032594599 -1882932396
      11'h6ba: T=64'b1100001010011111111100101101010110001111101011001001100010010000;  // -1029705003 -1884514160
      11'h6bb: T=64'b1100001011001100000100111100011110001111100101001000011100011110;  // -1026812985 -1886091490
      11'h6bc: T=64'b1100001011111000001111100010101110001111011111001000011100000010;  // -1023918549 -1887664382
      11'h6bd: T=64'b1100001100100100011100011111011110001111011001001001100001000000;  // -1021021705 -1889232832
      11'h6be: T=64'b1100001101010000101011110010011010001111010011001011101011011100;  // -1018122458 -1890796836
      11'h6bf: T=64'b1100001101111100111101011011000110001111001101001110111011011001;  // -1015220815 -1892356391
      11'h6c0: T=64'b1100001110101001010001011001000010001111000111010011010000111011;  // -1012316784 -1893911493
      11'h6c1: T=64'b1100001111010101100111101011111010001111000001011000101100000101;  // -1009410370 -1895462139
      11'h6c2: T=64'b1100010000000010000000010011001110001110111011011111001100111100;  // -1006501581 -1897008324
      11'h6c3: T=64'b1100010000101110011011001110100110001110110101100110110011100010;  // -1003590423 -1898550046
      11'h6c4: T=64'b1100010001011010111000011101011110001110101111101111011111111100;  // -1000676905 -1900087300
      11'h6c5: T=64'b1100010010000111010111111111100110001110101001111001010010001101;  // -997761031 -1901620083
      11'h6c6: T=64'b1100010010110011111001110100011110001110100100000100001010011001;  // -994842809 -1903148391
      11'h6c7: T=64'b1100010011100000011101111011100110001110011110010000001000100011;  // -991922247 -1904672221
      11'h6c8: T=64'b1100010100001101000100010100100110001110011000011101001100101111;  // -988999351 -1906191569
      11'h6c9: T=64'b1100010100111001101100111111000110001110010010101011010111000000;  // -986074127 -1907706432
      11'h6ca: T=64'b1100010101100110010111111010100110001110001100111010100111011010;  // -983146583 -1909216806
      11'h6cb: T=64'b1100010110010011000101000110101110001110000111001010111110000001;  // -980216725 -1910722687
      11'h6cc: T=64'b1100010110111111110100100010111110001110000001011100011010111000;  // -977284561 -1912224072
      11'h6cd: T=64'b1100010111101100100110001110111010001101111011101110111110000011;  // -974350098 -1913720957
      11'h6ce: T=64'b1100011000011001011010001010001110001101110110000010100111100101;  // -971413341 -1915213339
      11'h6cf: T=64'b1100011001000110010000010100010110001101110000010111010111100001;  // -968474299 -1916701215
      11'h6d0: T=64'b1100011001110011001000101100111010001101101010101101001101111100;  // -965532978 -1918184580
      11'h6d1: T=64'b1100011010100000000011010011011110001101100101000100001010111000;  // -962589385 -1919663432
      11'h6d2: T=64'b1100011011001101000000000111100110001101011111011100001110011010;  // -959643527 -1921137766
      11'h6d3: T=64'b1100011011111001111111001000111010001101011001110101011000100100;  // -956695410 -1922607580
      11'h6d4: T=64'b1100011100100111000000010110110110001101010100001111101001011010;  // -953745043 -1924072870
      11'h6d5: T=64'b1100011101010100000011110001000110001101001110101011000001000000;  // -950792431 -1925533632
      11'h6d6: T=64'b1100011110000001001001010111001010001101001001000111011111011001;  // -947837582 -1926989863
      11'h6d7: T=64'b1100011110101110010001001000101010001101000011100101000100101000;  // -944880502 -1928441560
      11'h6d8: T=64'b1100011111011011011011000101000010001100111110000011110000110001;  // -941921200 -1929888719
      11'h6d9: T=64'b1100100000001000100111001100000010001100111000100011100011110111;  // -938959680 -1931331337
      11'h6da: T=64'b1100100000110101110101011101000010001100110011000100011101111110;  // -935995952 -1932769410
      11'h6db: T=64'b1100100001100011000101110111110010001100101101100110011111001001;  // -933030020 -1934202935
      11'h6dc: T=64'b1100100010010000011000011011101010001100101000001001100111011011;  // -930061894 -1935631909
      11'h6dd: T=64'b1100100010111101101101001000011010001100100010101101110110111000;  // -927091578 -1937056328
      11'h6de: T=64'b1100100011101011000011111101011010001100011101010011001101100011;  // -924119082 -1938476189
      11'h6df: T=64'b1100100100011000011100111010011010001100010111111001101011011111;  // -921144410 -1939891489
      11'h6e0: T=64'b1100100101000101110111111110110110001100010010100001010000110000;  // -918167571 -1941302224
      11'h6e1: T=64'b1100100101110011010101001010010010001100001101001001111101011001;  // -915188572 -1942708391
      11'h6e2: T=64'b1100100110100000110100011100010110001100000111110011110001011110;  // -912207419 -1944109986
      11'h6e3: T=64'b1100100111001110010101110100100010001100000010011110101101000001;  // -909224120 -1945507007
      11'h6e4: T=64'b1100100111111011111001010010011110001011111101001010110000000110;  // -906238681 -1946899450
      11'h6e5: T=64'b1100101000101001011110110101101110001011110111110111111010110001;  // -903251109 -1948287311
      11'h6e6: T=64'b1100101001010111000110011101110010001011110010100110001101000100;  // -900261412 -1949670588
      11'h6e7: T=64'b1100101010000100110000001010001110001011101101010101100111000010;  // -897269597 -1951049278
      11'h6e8: T=64'b1100101010110010011011111010101010001011101000000110001000110000;  // -894275670 -1952423376
      11'h6e9: T=64'b1100101011100000001001101110100010001011100010110111110010010000;  // -891279640 -1953792880
      11'h6ea: T=64'b1100101100001101111001100101100110001011011101101010100011100101;  // -888281511 -1955157787
      11'h6eb: T=64'b1100101100111011101011011111001110001011011000011110011100110011;  // -885281293 -1956518093
      11'h6ec: T=64'b1100101101101001011111011011000110001011010011010011011101111101;  // -882278991 -1957873795
      11'h6ed: T=64'b1100101110010111010101011000101010001011001110001001100111000110;  // -879274614 -1959224890
      11'h6ee: T=64'b1100101111000101001101010111100110001011001001000000111000010010;  // -876268167 -1960571374
      11'h6ef: T=64'b1100101111110011000111010111011010001011000011111001010001100010;  // -873259658 -1961913246
      11'h6f0: T=64'b1100110000100001000011010111100110001010111110110010110010111100;  // -870249095 -1963250500
      11'h6f1: T=64'b1100110001001111000001010111110010001010111001101101011100100001;  // -867236484 -1964583135
      11'h6f2: T=64'b1100110001111101000001010111100010001010110100101001001110010101;  // -864221832 -1965911147
      11'h6f3: T=64'b1100110010101011000011010110011010001010101111100110001000011010;  // -861205146 -1967234534
      11'h6f4: T=64'b1100110011011001000111010011111010001010101010100100001010110101;  // -858186434 -1968553291
      11'h6f5: T=64'b1100110100000111001101001111100110001010100101100011010101101000;  // -855165703 -1969867416
      11'h6f6: T=64'b1100110100110101010101001001000110001010100000100011101000110111;  // -852142959 -1971176905
      11'h6f7: T=64'b1100110101100011011110111111111010001010011011100101000100100100;  // -849118210 -1972481756
      11'h6f8: T=64'b1100110110010001101010110011100110001010010110100111101000110010;  // -846091463 -1973781966
      11'h6f9: T=64'b1100110110111111111000100011101110001010010001101011010101100100;  // -843062725 -1975077532
      11'h6fa: T=64'b1100110111101110001000001111110110001010001100110000001010111111;  // -840032003 -1976368449
      11'h6fb: T=64'b1100111000011100011001110111011110001010000111110110001001000100;  // -836999305 -1977654716
      11'h6fc: T=64'b1100111001001010101101011010001110001010000010111101001111110110;  // -833964637 -1978936330
      11'h6fd: T=64'b1100111001111001000010110111100110001001111110000101011111011001;  // -830928007 -1980213287
      11'h6fe: T=64'b1100111010100111011010001111001110001001111001001110110111110000;  // -827889421 -1981485584
      11'h6ff: T=64'b1100111011010101110011100000100010001001110100011001011000111101;  // -824848888 -1982753219
      11'h700: T=64'b1100111100000100001110101011001110001001101111100101000011000100;  // -821806413 -1984016188
      11'h701: T=64'b1100111100110010101011101110101110001001101010110001110110001000;  // -818762005 -1985274488
      11'h702: T=64'b1100111101100001001010101010101010001001100101111111110010001011;  // -815715670 -1986528117
      11'h703: T=64'b1100111110001111101011011110100110001001100001001110110111010000;  // -812667415 -1987777072
      11'h704: T=64'b1100111110111110001110001010000010001001011100011111000101011011;  // -809617248 -1989021349
      11'h705: T=64'b1100111111101100110010101100100010001001010111110000011100101111;  // -806565176 -1990260945
      11'h706: T=64'b1101000000011011011001000101100110001001010011000010111101001101;  // -803511207 -1991495859
      11'h707: T=64'b1101000001001010000001010100111010001001001110010110100110111010;  // -800455346 -1992726086
      11'h708: T=64'b1101000001111000101011011001111010001001001001101011011001111000;  // -797397602 -1993951624
      11'h709: T=64'b1101000010100111010111010100001110001001000101000001010110001010;  // -794337981 -1995172470
      11'h70a: T=64'b1101000011010110000101000011010010001001000000011000011011110011;  // -791276492 -1996388621
      11'h70b: T=64'b1101000100000100110100100110110010001000111011110000101010110101;  // -788213140 -1997600075
      11'h70c: T=64'b1101000100110011100101111110001010001000110111001010000011010100;  // -785147934 -1998806828
      11'h70d: T=64'b1101000101100010011001001001000010001000110010100100100101010010;  // -782080880 -2000008878
      11'h70e: T=64'b1101000110010001001110000110111010001000101110000000010000110011;  // -779011986 -2001206221
      11'h70f: T=64'b1101000111000000000100110111010110001000101001011101000101111000;  // -775941259 -2002398856
      11'h710: T=64'b1101000111101110111101011001111010001000100100111011000100100110;  // -772868706 -2003586778
      11'h711: T=64'b1101001000011101110111101110001010001000100000011010001100111110;  // -769794334 -2004769986
      11'h712: T=64'b1101001001001100110011110011100110001000011011111010011111000011;  // -766718151 -2005948477
      11'h713: T=64'b1101001001111011110001101001110110001000010111011011111010111001;  // -763640163 -2007122247
      11'h714: T=64'b1101001010101010110001010000010110001000010010111110100000100001;  // -760560379 -2008291295
      11'h715: T=64'b1101001011011001110010100110101110001000001110100010010000000000;  // -757478805 -2009455616
      11'h716: T=64'b1101001100001000110101101100011110001000001010000111001001010111;  // -754395449 -2010615209
      11'h717: T=64'b1101001100110111111010100001001010001000000101101101001100101000;  // -751310318 -2011770072
      11'h718: T=64'b1101001101100111000001000100011010001000000001010100011001111000;  // -748223418 -2012920200
      11'h719: T=64'b1101001110010110001001010101101010000111111100111100110001001001;  // -745134758 -2014065591
      11'h71a: T=64'b1101001111000101010011010100011110000111111000100110010010011100;  // -742044345 -2015206244
      11'h71b: T=64'b1101001111110100011111000000011110000111110100010000111101110110;  // -738952185 -2016342154
      11'h71c: T=64'b1101010000100011101100011001000110000111101111111100110011011000;  // -735858287 -2017473320
      11'h71d: T=64'b1101010001010010111011011101111110000111101011101001110011000110;  // -732762657 -2018599738
      11'h71e: T=64'b1101010010000010001100001110100110000111100111010111111101000001;  // -729665303 -2019721407
      11'h71f: T=64'b1101010010110001011110101010100010000111100011000111010001001110;  // -726566232 -2020838322
      11'h720: T=64'b1101010011100000110010110001010110000111011110110111101111101101;  // -723465451 -2021950483
      11'h721: T=64'b1101010100010000001000100010100010000111011010101001011000100010;  // -720362968 -2023057886
      11'h722: T=64'b1101010100111111011111111101101010000111010110011100001011110000;  // -717258790 -2024160528
      11'h723: T=64'b1101010101101110111001000010010010000111010010010000001001011001;  // -714152924 -2025258407
      11'h724: T=64'b1101010110011110010011101111111110000111001110000101010001011111;  // -711045377 -2026351521
      11'h725: T=64'b1101010111001101110000000110001110000111001001111011100100000110;  // -707936157 -2027439866
      11'h726: T=64'b1101010111111101001110000100100010000111000101110011000001001111;  // -704825272 -2028523441
      11'h727: T=64'b1101011000101100101101101010100010000111000001101011101000111110;  // -701712728 -2029602242
      11'h728: T=64'b1101011001011100001110110111101110000110111101100101011011010100;  // -698598533 -2030676268
      11'h729: T=64'b1101011010001011110001101011101010000110111001100000011000010101;  // -695482694 -2031745515
      11'h72a: T=64'b1101011010111011010110000101111010000110110101011100100000000011;  // -692365218 -2032809981
      11'h72b: T=64'b1101011011101010111100000101111110000110110001011001110010100000;  // -689246113 -2033869664
      11'h72c: T=64'b1101011100011010100011101011011010000110101101011000001111101111;  // -686125386 -2034924561
      11'h72d: T=64'b1101011101001010001100110101101110000110101001010111110111110011;  // -683003045 -2035974669
      11'h72e: T=64'b1101011101111001110111100100011110000110100101011000101010101101;  // -679879097 -2037019987
      11'h72f: T=64'b1101011110101001100011110111001110000110100001011010101000100000;  // -676753549 -2038060512
      11'h730: T=64'b1101011111011001010001101101100010000110011101011101110001010000;  // -673626408 -2039096240
      11'h731: T=64'b1101100000001001000001000110111010000110011001100010000100111101;  // -670497682 -2040127171
      11'h732: T=64'b1101100000111000110010000010110110000110010101100111100011101011;  // -667367379 -2041153301
      11'h733: T=64'b1101100001101000100100100000111110000110010001101110001101011101;  // -664235505 -2042174627
      11'h734: T=64'b1101100010011000011000100000110010000110001101110110000010010011;  // -661102068 -2043191149
      11'h735: T=64'b1101100011001000001110000001110110000110001001111111000010010010;  // -657967075 -2044202862
      11'h736: T=64'b1101100011111000000101000011101010000110000110001001001101011010;  // -654830534 -2045209766
      11'h737: T=64'b1101100100100111111101100101101110000110000010010100100011110000;  // -651692453 -2046211856
      11'h738: T=64'b1101100101010111110111100111101110000101111110100001000101010100;  // -648552837 -2047209132
      11'h739: T=64'b1101100110000111110011001001000010000101111010101110110010001001;  // -645411696 -2048201591
      11'h73a: T=64'b1101100110110111110000001001010010000101110110111101101010010010;  // -642269036 -2049189230
      11'h73b: T=64'b1101100111100111101110100111111110000101110011001101101101110001;  // -639124865 -2050172047
      11'h73c: T=64'b1101101000010111101110100100101010000101101111011110111100101000;  // -635979190 -2051150040
      11'h73d: T=64'b1101101001000111101111111110111010000101101011110001010110111010;  // -632832018 -2052123206
      11'h73e: T=64'b1101101001110111110010110110001110000101101000000100111100101001;  // -629683357 -2053091543
      11'h73f: T=64'b1101101010100111110111001010001010000101100100011001101101110111;  // -626533214 -2054055049
      11'h740: T=64'b1101101011010111111100111010001110000101100000101111101010100110;  // -623381597 -2055013722
      11'h741: T=64'b1101101100001000000100000101111010000101011101000110110010111001;  // -620228514 -2055967559
      11'h742: T=64'b1101101100111000001100101100111010000101011001011111000110110001;  // -617073970 -2056916559
      11'h743: T=64'b1101101101101000010110101110100110000101010101111000100110010010;  // -613917975 -2057860718
      11'h744: T=64'b1101101110011000100010001010100110000101010010010011010001011101;  // -610760535 -2058800035
      11'h745: T=64'b1101101111001000101111000000011010000101001110101111001000010101;  // -607601658 -2059734507
      11'h746: T=64'b1101101111111000111101001111100110000101001011001100001010111100;  // -604441351 -2060664132
      11'h747: T=64'b1101110000101001001100110111101010000101000111101010011001010011;  // -601279622 -2061588909
      11'h748: T=64'b1101110001011001011101111000001010000101000100001001110011011101;  // -598116478 -2062508835
      11'h749: T=64'b1101110010001001110000010000100110000101000000101010011001011101;  // -594951927 -2063423907
      11'h74a: T=64'b1101110010111010000100000000100010000100111101001100001011010101;  // -591785976 -2064334123
      11'h74b: T=64'b1101110011101010011001000111100010000100111001101111001001000101;  // -588618632 -2065239483
      11'h74c: T=64'b1101110100011010101111100101000110000100110110010011010010110010;  // -585449903 -2066139982
      11'h74d: T=64'b1101110101001011000111011000110010000100110010111000101000011100;  // -582279796 -2067035620
      11'h74e: T=64'b1101110101111011100000100010000110000100101111011111001010000111;  // -579108319 -2067926393
      11'h74f: T=64'b1101110110101011111011000000100010000100101100000110110111110011;  // -575935480 -2068812301
      11'h750: T=64'b1101110111011100010110110011101110000100101000101111110001100011;  // -572761285 -2069693341
      11'h751: T=64'b1101111000001100110011111011000110000100100101011001110111011010;  // -569585743 -2070569510
      11'h752: T=64'b1101111000111101010010010110010010000100100010000101001001011001;  // -566408860 -2071440807
      11'h753: T=64'b1101111001101101110010000100110010000100011110110001100111100010;  // -563230644 -2072307230
      11'h754: T=64'b1101111010011110010011000110000110000100011011011111010001111000;  // -560051103 -2073168776
      11'h755: T=64'b1101111011001110110101011001101110000100011000001110001000011011;  // -556870245 -2074025445
      11'h756: T=64'b1101111011111111011000111111010010000100010100111110001011010000;  // -553688076 -2074877232
      11'h757: T=64'b1101111100101111111101110110010010000100010001101111011010010110;  // -550504604 -2075724138
      11'h758: T=64'b1101111101100000100011111110010010000100001110100001110101110001;  // -547319836 -2076566159
      11'h759: T=64'b1101111110010001001011010110101110000100001011010101011101100011;  // -544133781 -2077403293
      11'h75a: T=64'b1101111111000001110011111111001110000100001000001010010001101101;  // -540946445 -2078235539
      11'h75b: T=64'b1101111111110010011101110111001110000100000101000000010010010001;  // -537757837 -2079062895
      11'h75c: T=64'b1110000000100011001000111110010110000100000001110111011111010001;  // -534567963 -2079885359
      11'h75d: T=64'b1110000001010011110101010100000110000011111110101111111000101111;  // -531376831 -2080702929
      11'h75e: T=64'b1110000010000100100010111000000010000011111011101001011110101110;  // -528184448 -2081515602
      11'h75f: T=64'b1110000010110101010001101001100110000011111000100100010001001110;  // -524990823 -2082323378
      11'h760: T=64'b1110000011100110000001101000010110000011110101100000010000010011;  // -521795963 -2083126253
      11'h761: T=64'b1110000100010110110010110011110110000011110010011101011011111101;  // -518599875 -2083924227
      11'h762: T=64'b1110000101000111100101001011101010000011101111011011110100001111;  // -515402566 -2084717297
      11'h763: T=64'b1110000101111000011000101111001110000011101100011011011001001010;  // -512204045 -2085505462
      11'h764: T=64'b1110000110101001001101011110001010000011101001011100001010110001;  // -509004318 -2086288719
      11'h765: T=64'b1110000111011010000011010111111110000011100110011110001001000101;  // -505803393 -2087067067
      11'h766: T=64'b1110001000001010111010011100000110000011100011100001010100001000;  // -502601279 -2087840504
      11'h767: T=64'b1110001000111011110010101010001110000011100000100101101011111100;  // -499397981 -2088609028
      11'h768: T=64'b1110001001101100101100000001101110000011011101101011010000100011;  // -496193509 -2089372637
      11'h769: T=64'b1110001010011101100110100010001110000011011010110010000001111110;  // -492987869 -2090131330
      11'h76a: T=64'b1110001011001110100010001011001110000011010111111010000000010000;  // -489781069 -2090885104
      11'h76b: T=64'b1110001011111111011110111100010010000011010101000011001011011001;  // -486573116 -2091633959
      11'h76c: T=64'b1110001100110000011100110100110110000011010010001101100011011101;  // -483364019 -2092377891
      11'h76d: T=64'b1110001101100001011011110100100010000011001111011001001000011100;  // -480153784 -2093116900
      11'h76e: T=64'b1110001110010010011011111010110110000011001100100101111010011000;  // -476942419 -2093850984
      11'h76f: T=64'b1110001111000011011101000111010010000011001001110011111001010011;  // -473729932 -2094580141
      11'h770: T=64'b1110001111110100011111011001011010000011000111000011000101001111;  // -470516330 -2095304369
      11'h771: T=64'b1110010000100101100010110000101110000011000100010011011110001110;  // -467301621 -2096023666
      11'h772: T=64'b1110010001010110100111001100101110000011000001100101000100010001;  // -464085813 -2096738031
      11'h773: T=64'b1110010010000111101100101101000010000010111110110111110111011001;  // -460868912 -2097447463
      11'h774: T=64'b1110010010111000110011010001000110000010111100001011110111101001;  // -457650927 -2098151959
      11'h775: T=64'b1110010011101001111010111000011110000010111001100001000101000010;  // -454431865 -2098851518
      11'h776: T=64'b1110010100011011000011100010101010000010110110110111011111100110;  // -451211734 -2099546138
      11'h777: T=64'b1110010101001100001101001111001110000010110100001111000111010110;  // -447990541 -2100235818
      11'h778: T=64'b1110010101111101010111111101101110000010110001100111111100010101;  // -444768293 -2100920555
      11'h779: T=64'b1110010110101110100011101101100010000010101111000001111110100011;  // -441545000 -2101600349
      11'h77a: T=64'b1110010111011111110000011110010110000010101100011101001110000010;  // -438320667 -2102275198
      11'h77b: T=64'b1110011000010000111110001111100110000010101001111001101010110100;  // -435095303 -2102945100
      11'h77c: T=64'b1110011001000010001101000000110110000010100111010111010100111011;  // -431868915 -2103610053
      11'h77d: T=64'b1110011001110011011100110001101010000010100100110110001100011000;  // -428641510 -2104270056
      11'h77e: T=64'b1110011010100100101101100001011010000010100010010110010001001100;  // -425413098 -2104925108
      11'h77f: T=64'b1110011011010101111111001111110010000010011111110111100011011001;  // -422183684 -2105575207
      11'h780: T=64'b1110011100000111010001111100010010000010011101011010000011000001;  // -418953276 -2106220351
      11'h781: T=64'b1110011100111000100101100110010110000010011010111101110000000101;  // -415721883 -2106860539
      11'h782: T=64'b1110011101101001111010001101100010000010011000100010101010100111;  // -412489512 -2107495769
      11'h783: T=64'b1110011110011011001111110001011010000010010110001000110010101000;  // -409256170 -2108126040
      11'h784: T=64'b1110011111001100100110010001100010000010010011110000001000001001;  // -406021864 -2108751351
      11'h785: T=64'b1110011111111101111101101101010010000010010001011000101011001101;  // -402786604 -2109371699
      11'h786: T=64'b1110100000101111010110000100010010000010001111000010011011110100;  // -399550396 -2109987084
      11'h787: T=64'b1110100001100000101111010110000110000010001100101101011010000000;  // -396313247 -2110597504
      11'h788: T=64'b1110100010010010001001100010001010000010001010011001100101110010;  // -393075166 -2111202958
      11'h789: T=64'b1110100011000011100100101000000010000010001000000110111111001101;  // -389836160 -2111803443
      11'h78a: T=64'b1110100011110101000000100111001110000010000101110101100110010001;  // -386596237 -2112398959
      11'h78b: T=64'b1110100100100110011101011111010010000010000011100101011010111111;  // -383355404 -2112989505
      11'h78c: T=64'b1110100101010111111011001111101110000010000001010110011101011001;  // -380113669 -2113575079
      11'h78d: T=64'b1110100110001001011001111000000110000001111111001000101101100001;  // -376871039 -2114155679
      11'h78e: T=64'b1110100110111010111001010111110110000001111100111100001011011000;  // -373627523 -2114731304
      11'h78f: T=64'b1110100111101100011001101110100110000001111010110000110110111111;  // -370383127 -2115301953
      11'h790: T=64'b1110101000011101111010111011110010000001111000100110110000010111;  // -367137860 -2115867625
      11'h791: T=64'b1110101001001111011100111110111110000001110110011101110111100010;  // -363891729 -2116428318
      11'h792: T=64'b1110101010000000111111110111101010000001110100010110001100100010;  // -360644742 -2116984030
      11'h793: T=64'b1110101010110010100011100101011010000001110010001111101111010111;  // -357396906 -2117534761
      11'h794: T=64'b1110101011100100001000000111101110000001110000001010100000000010;  // -354148229 -2118080510
      11'h795: T=64'b1110101100010101101101011110000110000001101110000110011110100110;  // -350898719 -2118621274
      11'h796: T=64'b1110101101000111010011101000000110000001101100000011101011000011;  // -347648383 -2119157053
      11'h797: T=64'b1110101101111000111010100101001110000001101010000010000101011010;  // -344397229 -2119687846
      11'h798: T=64'b1110101110101010100010010100111110000001101000000001101101101110;  // -341145265 -2120213650
      11'h799: T=64'b1110101111011100001010110110111010000001100110000010100011111110;  // -337892498 -2120734466
      11'h79a: T=64'b1110110000001101110100001010100010000001100100000100101000001101;  // -334638936 -2121250291
      11'h79b: T=64'b1110110000111111011110001111011010000001100010000111111010011011;  // -331384586 -2121761125
      11'h79c: T=64'b1110110001110001001001000100111110000001100000001100011010101010;  // -328129457 -2122266966
      11'h79d: T=64'b1110110010100010110100101010110110000001011110010010001000111011;  // -324873555 -2122767813
      11'h79e: T=64'b1110110011010100100001000000011110000001011100011001000101001111;  // -321616889 -2123263665
      11'h79f: T=64'b1110110100000110001110000101011010000001011010100001001111100111;  // -318359466 -2123754521
      11'h7a0: T=64'b1110110100110111111011111001001010000001011000101010101000000101;  // -315101294 -2124240379
      11'h7a1: T=64'b1110110101101001101010011011001110000001010110110101001110101001;  // -311842381 -2124721239
      11'h7a2: T=64'b1110110110011011011001101011001010000001010101000001000011010101;  // -308582734 -2125197099
      11'h7a3: T=64'b1110110111001101001001101000011110000001010011001110000110001001;  // -305322361 -2125667959
      11'h7a4: T=64'b1110110111111110111010010010101110000001010001011100010111001000;  // -302061269 -2126133816
      11'h7a5: T=64'b1110111000110000101011101001011010000001001111101011110110010001;  // -298799466 -2126594671
      11'h7a6: T=64'b1110111001100010011101101011111110000001001101111100100011100111;  // -295536961 -2127050521
      11'h7a7: T=64'b1110111010010100010000011010000010000001001100001110011111001010;  // -292273760 -2127501366
      11'h7a8: T=64'b1110111011000110000011110011000110000001001010100001101000111011;  // -289009871 -2127947205
      11'h7a9: T=64'b1110111011110111110111110110101010000001001000110110000000111011;  // -285745302 -2128388037
      11'h7aa: T=64'b1110111100101001101100100100001110000001000111001011100111001011;  // -282480061 -2128823861
      11'h7ab: T=64'b1110111101011011100001111011010110000001000101100010011011101101;  // -279214155 -2129254675
      11'h7ac: T=64'b1110111110001101010111111011100010000001000011111010011110100001;  // -275947592 -2129680479
      11'h7ad: T=64'b1110111110111111001110100100010110000001000010010011101111101001;  // -272680379 -2130101271
      11'h7ae: T=64'b1110111111110001000101110101001110000001000000101110001111000101;  // -269412525 -2130517051
      11'h7af: T=64'b1111000000100010111101101101101110000000111111001001111100110110;  // -266144037 -2130927818
      11'h7b0: T=64'b1111000001010100110110001101010110000000111101100110111000111101;  // -262874923 -2131333571
      11'h7b1: T=64'b1111000010000110101111010011101010000000111100000101000011011100;  // -259605190 -2131734308
      11'h7b2: T=64'b1111000010111000101001000000000110000000111010100100011100010011;  // -256334847 -2132130029
      11'h7b3: T=64'b1111000011101010100011010010010010000000111001000101000011100011;  // -253063900 -2132520733
      11'h7b4: T=64'b1111000100011100011110001001101010000000110111100110111001001101;  // -249792358 -2132906419
      11'h7b5: T=64'b1111000101001110011001100101110010000000110110001001111101010010;  // -246520228 -2133287086
      11'h7b6: T=64'b1111000110000000010101100110001110000000110100101110001111110011;  // -243247517 -2133662733
      11'h7b7: T=64'b1111000110110010010010001010010110000000110011010011110000110000;  // -239974235 -2134033360
      11'h7b8: T=64'b1111000111100100001111010001110010000000110001111010100000001011;  // -236700388 -2134398965
      11'h7b9: T=64'b1111001000010110001100111100000110000000110000100010011110000101;  // -233425983 -2134759547
      11'h7ba: T=64'b1111001001001000001011001000101010000000101111001011101010011110;  // -230151030 -2135115106
      11'h7bb: T=64'b1111001001111010001001110111000110000000101101110110000101010111;  // -226875535 -2135465641
      11'h7bc: T=64'b1111001010101100001001000110111010000000101100100001101110110000;  // -223599506 -2135811152
      11'h7bd: T=64'b1111001011011110001000110111100110000000101011001110100110101100;  // -220322951 -2136151636
      11'h7be: T=64'b1111001100010000001001001000101110000000101001111100101101001010;  // -217045877 -2136487094
      11'h7bf: T=64'b1111001101000010001001111001101110000000101000101100000010001100;  // -213768293 -2136817524
      11'h7c0: T=64'b1111001101110100001011001010001010000000100111011100100101110010;  // -210490206 -2137142926
      11'h7c1: T=64'b1111001110100110001100111001100110000000100110001110010111111100;  // -207211623 -2137463300
      11'h7c2: T=64'b1111001111011000001111000111011110000000100101000001011000101101;  // -203932553 -2137778643
      11'h7c3: T=64'b1111010000001010010001110011010110000000100011110101101000000011;  // -200653003 -2138088957
      11'h7c4: T=64'b1111010000111100010100111100101110000000100010101011000110000001;  // -197372981 -2138394239
      11'h7c5: T=64'b1111010001101110011000100011001010000000100001100001110010100111;  // -194092494 -2138694489
      11'h7c6: T=64'b1111010010100000011100100110000110000000100000011001101101110101;  // -190811551 -2138989707
      11'h7c7: T=64'b1111010011010010100001000101000110000000011111010010110111101101;  // -187530159 -2139279891
      11'h7c8: T=64'b1111010100000100100101111111101110000000011110001101010000001110;  // -184248325 -2139565042
      11'h7c9: T=64'b1111010100110110101011010101011010000000011101001000110111011010;  // -180966058 -2139845158
      11'h7ca: T=64'b1111010101101000110001000101101110000000011100000101101101010001;  // -177683365 -2140120239
      11'h7cb: T=64'b1111010110011010110111010000001010000000011011000011110001110101;  // -174400254 -2140390283
      11'h7cc: T=64'b1111010111001100111101110100010010000000011010000011000101000100;  // -171116732 -2140655292
      11'h7cd: T=64'b1111010111111111000100110001100010000000011001000011100111000001;  // -167832808 -2140915263
      11'h7ce: T=64'b1111011000110001001100000111011110000000011000000101010111101100;  // -164548489 -2141170196
      11'h7cf: T=64'b1111011001100011010011110101100110000000010111001000010111000101;  // -161263783 -2141420091
      11'h7d0: T=64'b1111011010010101011011111011011110000000010110001100100101001101;  // -157978697 -2141664947
      11'h7d1: T=64'b1111011011000111100100011000100010000000010101010010000010000101;  // -154693240 -2141904763
      11'h7d2: T=64'b1111011011111001101101001100011010000000010100011000101101101100;  // -151407418 -2142139540
      11'h7d3: T=64'b1111011100101011110110010110011110000000010011100000101000000101;  // -148121241 -2142369275
      11'h7d4: T=64'b1111011101011101111111110110011010000000010010101001110001001110;  // -144834714 -2142593970
      11'h7d5: T=64'b1111011110010000001001101011100110000000010001110100001001001001;  // -141547847 -2142813623
      11'h7d6: T=64'b1111011111000010010011110101100110000000010000111111101111110111;  // -138260647 -2143028233
      11'h7d7: T=64'b1111011111110100011110010011111010000000010000001100100101010111;  // -134973122 -2143237801
      11'h7d8: T=64'b1111100000100110101001000110001010000000001111011010101001101011;  // -131685278 -2143442325
      11'h7d9: T=64'b1111100001011000110100001011101110000000001110101001111100110010;  // -128397125 -2143641806
      11'h7da: T=64'b1111100010001010111111100100001010000000001101111010011110101101;  // -125108670 -2143836243
      11'h7db: T=64'b1111100010111101001011001110111110000000001101001100001111011110;  // -121819921 -2144025634
      11'h7dc: T=64'b1111100011101111010111001011101110000000001100011111001111000011;  // -118530885 -2144209981
      11'h7dd: T=64'b1111100100100001100011011001111010000000001011110011011101011110;  // -115241570 -2144389282
      11'h7de: T=64'b1111100101010011101111111001000110000000001011001000111010101110;  // -111951983 -2144563538
      11'h7df: T=64'b1111100110000101111100101000101010000000001010011111100110110101;  // -108662134 -2144732747
      11'h7e0: T=64'b1111100110111000001001101000010010000000001001110111100001110011;  // -105372028 -2144896909
      11'h7e1: T=64'b1111100111101010010110110111010110000000001001010000101011101000;  // -102081675 -2145056024
      11'h7e2: T=64'b1111101000011100100100010101011110000000001000101011000100010101;  // -98791081 -2145210091
      11'h7e3: T=64'b1111101001001110110010000010000110000000001000000110101011111001;  // -95500255 -2145359111
      11'h7e4: T=64'b1111101010000000111111111100101110000000000111100011100010010110;  // -92209205 -2145503082
      11'h7e5: T=64'b1111101010110011001110000100111110000000000111000001100111101011;  // -88917937 -2145642005
      11'h7e6: T=64'b1111101011100101011100011010010010000000000110100000111011111001;  // -85626460 -2145775879
      11'h7e7: T=64'b1111101100010111101010111100001010000000000110000001011111000000;  // -82334782 -2145904704
      11'h7e8: T=64'b1111101101001001111001101010001110000000000101100011010001000001;  // -79042909 -2146028479
      11'h7e9: T=64'b1111101101111100001000100011110110000000000101000110010001111100;  // -75750851 -2146147204
      11'h7ea: T=64'b1111101110101110010111101000100110000000000100101010100001110000;  // -72458615 -2146260880
      11'h7eb: T=64'b1111101111100000100110111000000010000000000100010000000000100000;  // -69166208 -2146369504
      11'h7ec: T=64'b1111110000010010110110010001101010000000000011110110101110001001;  // -65873638 -2146473079
      11'h7ed: T=64'b1111110001000101000101110100111010000000000011011110101010101110;  // -62580914 -2146571602
      11'h7ee: T=64'b1111110001110111010101100001011010000000000011000111110110001101;  // -59288042 -2146665075
      11'h7ef: T=64'b1111110010101001100101010110101010000000000010110010010000101000;  // -55995030 -2146753496
      11'h7f0: T=64'b1111110011011011110101010100000110000000000010011101111001111111;  // -52701887 -2146836865
      11'h7f1: T=64'b1111110100001110000101011001010010000000000010001010110010010001;  // -49408620 -2146915183
      11'h7f2: T=64'b1111110101000000010101100101110010000000000001111000111001011111;  // -46115236 -2146988449
      11'h7f3: T=64'b1111110101110010100101111001000010000000000001101000001111101001;  // -42821744 -2147056663
      11'h7f4: T=64'b1111110110100100110110010010100110000000000001011000110100110000;  // -39528151 -2147119824
      11'h7f5: T=64'b1111110111010111000110110001111010000000000001001010101000110011;  // -36234466 -2147177933
      11'h7f6: T=64'b1111111000001001010111010110100110000000000000111101101011110010;  // -32940695 -2147230990
      11'h7f7: T=64'b1111111000111011101000000000001010000000000000110001111101101110;  // -29646846 -2147278994
      11'h7f8: T=64'b1111111001101101111000101110000010000000000000100111011110100111;  // -26352928 -2147321945
      11'h7f9: T=64'b1111111010100000001001011111110110000000000000011110001110011100;  // -23058947 -2147359844
      11'h7fa: T=64'b1111111011010010011010010100111110000000000000010110001101001111;  // -19764913 -2147392689
      11'h7fb: T=64'b1111111100000100101011001101000010000000000000001111011010111110;  // -16470832 -2147420482
      11'h7fc: T=64'b1111111100110110111100000111100010000000000000001001110111101011;  // -13176712 -2147443221
      11'h7fd: T=64'b1111111101101001001101000011111110000000000000000101100011010101;  // -9882561 -2147460907
      11'h7fe: T=64'b1111111110011011011110000001110110000000000000000010011101111011;  // -6588387 -2147473541
      11'h7ff: T=64'b1111111111001101101111000000101110000000000000000000100111100000;  // -3294197 -2147481120
      default: T=64'b0;
    endcase

endmodule
