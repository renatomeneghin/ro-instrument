`timescale 1ns/10ps

module COREDDS_C0_COREDDS_C0_0_dds_qrtr_cos (index, cosine);
  input  [8:0] index;
  output [17:0] cosine;
  reg signed [17:0] cosine/* synthesis syn_maxfan = 1000 */;

  always @ (index) 
    case (index) 
         0: cosine = 18'b010000000000000000;  //      65536 
         1: cosine = 18'b010000000000000000;  //      65536 
         2: cosine = 18'b010000000000000000;  //      65536 
         3: cosine = 18'b001111111111111111;  //      65535 
         4: cosine = 18'b001111111111111110;  //      65534 
         5: cosine = 18'b001111111111111110;  //      65534 
         6: cosine = 18'b001111111111111101;  //      65533 
         7: cosine = 18'b001111111111111100;  //      65532 
         8: cosine = 18'b001111111111111010;  //      65530 
         9: cosine = 18'b001111111111111001;  //      65529 
        10: cosine = 18'b001111111111110111;  //      65527 
        11: cosine = 18'b001111111111110110;  //      65526 
        12: cosine = 18'b001111111111110100;  //      65524 
        13: cosine = 18'b001111111111110010;  //      65522 
        14: cosine = 18'b001111111111110000;  //      65520 
        15: cosine = 18'b001111111111101101;  //      65517 
        16: cosine = 18'b001111111111101011;  //      65515 
        17: cosine = 18'b001111111111101000;  //      65512 
        18: cosine = 18'b001111111111100110;  //      65510 
        19: cosine = 18'b001111111111100011;  //      65507 
        20: cosine = 18'b001111111111100000;  //      65504 
        21: cosine = 18'b001111111111011100;  //      65500 
        22: cosine = 18'b001111111111011001;  //      65497 
        23: cosine = 18'b001111111111010101;  //      65493 
        24: cosine = 18'b001111111111010010;  //      65490 
        25: cosine = 18'b001111111111001110;  //      65486 
        26: cosine = 18'b001111111111001010;  //      65482 
        27: cosine = 18'b001111111111000110;  //      65478 
        28: cosine = 18'b001111111111000001;  //      65473 
        29: cosine = 18'b001111111110111101;  //      65469 
        30: cosine = 18'b001111111110111000;  //      65464 
        31: cosine = 18'b001111111110110100;  //      65460 
        32: cosine = 18'b001111111110101111;  //      65455 
        33: cosine = 18'b001111111110101001;  //      65449 
        34: cosine = 18'b001111111110100100;  //      65444 
        35: cosine = 18'b001111111110011111;  //      65439 
        36: cosine = 18'b001111111110011001;  //      65433 
        37: cosine = 18'b001111111110010100;  //      65428 
        38: cosine = 18'b001111111110001110;  //      65422 
        39: cosine = 18'b001111111110001000;  //      65416 
        40: cosine = 18'b001111111110000010;  //      65410 
        41: cosine = 18'b001111111101111011;  //      65403 
        42: cosine = 18'b001111111101110101;  //      65397 
        43: cosine = 18'b001111111101101110;  //      65390 
        44: cosine = 18'b001111111101100111;  //      65383 
        45: cosine = 18'b001111111101100000;  //      65376 
        46: cosine = 18'b001111111101011001;  //      65369 
        47: cosine = 18'b001111111101010010;  //      65362 
        48: cosine = 18'b001111111101001011;  //      65355 
        49: cosine = 18'b001111111101000011;  //      65347 
        50: cosine = 18'b001111111100111011;  //      65339 
        51: cosine = 18'b001111111100110100;  //      65332 
        52: cosine = 18'b001111111100101100;  //      65324 
        53: cosine = 18'b001111111100100011;  //      65315 
        54: cosine = 18'b001111111100011011;  //      65307 
        55: cosine = 18'b001111111100010011;  //      65299 
        56: cosine = 18'b001111111100001010;  //      65290 
        57: cosine = 18'b001111111100000001;  //      65281 
        58: cosine = 18'b001111111011111000;  //      65272 
        59: cosine = 18'b001111111011101111;  //      65263 
        60: cosine = 18'b001111111011100110;  //      65254 
        61: cosine = 18'b001111111011011101;  //      65245 
        62: cosine = 18'b001111111011010011;  //      65235 
        63: cosine = 18'b001111111011001001;  //      65225 
        64: cosine = 18'b001111111010111111;  //      65215 
        65: cosine = 18'b001111111010110101;  //      65205 
        66: cosine = 18'b001111111010101011;  //      65195 
        67: cosine = 18'b001111111010100001;  //      65185 
        68: cosine = 18'b001111111010010111;  //      65175 
        69: cosine = 18'b001111111010001100;  //      65164 
        70: cosine = 18'b001111111010000001;  //      65153 
        71: cosine = 18'b001111111001110110;  //      65142 
        72: cosine = 18'b001111111001101011;  //      65131 
        73: cosine = 18'b001111111001100000;  //      65120 
        74: cosine = 18'b001111111001010101;  //      65109 
        75: cosine = 18'b001111111001001001;  //      65097 
        76: cosine = 18'b001111111000111101;  //      65085 
        77: cosine = 18'b001111111000110001;  //      65073 
        78: cosine = 18'b001111111000100101;  //      65061 
        79: cosine = 18'b001111111000011001;  //      65049 
        80: cosine = 18'b001111111000001101;  //      65037 
        81: cosine = 18'b001111111000000001;  //      65025 
        82: cosine = 18'b001111110111110100;  //      65012 
        83: cosine = 18'b001111110111100111;  //      64999 
        84: cosine = 18'b001111110111011010;  //      64986 
        85: cosine = 18'b001111110111001101;  //      64973 
        86: cosine = 18'b001111110111000000;  //      64960 
        87: cosine = 18'b001111110110110011;  //      64947 
        88: cosine = 18'b001111110110100101;  //      64933 
        89: cosine = 18'b001111110110010111;  //      64919 
        90: cosine = 18'b001111110110001001;  //      64905 
        91: cosine = 18'b001111110101111100;  //      64892 
        92: cosine = 18'b001111110101101101;  //      64877 
        93: cosine = 18'b001111110101011111;  //      64863 
        94: cosine = 18'b001111110101010001;  //      64849 
        95: cosine = 18'b001111110101000010;  //      64834 
        96: cosine = 18'b001111110100110011;  //      64819 
        97: cosine = 18'b001111110100100100;  //      64804 
        98: cosine = 18'b001111110100010101;  //      64789 
        99: cosine = 18'b001111110100000110;  //      64774 
       100: cosine = 18'b001111110011110111;  //      64759 
       101: cosine = 18'b001111110011100111;  //      64743 
       102: cosine = 18'b001111110011011000;  //      64728 
       103: cosine = 18'b001111110011001000;  //      64712 
       104: cosine = 18'b001111110010111000;  //      64696 
       105: cosine = 18'b001111110010101000;  //      64680 
       106: cosine = 18'b001111110010010111;  //      64663 
       107: cosine = 18'b001111110010000111;  //      64647 
       108: cosine = 18'b001111110001110110;  //      64630 
       109: cosine = 18'b001111110001100110;  //      64614 
       110: cosine = 18'b001111110001010101;  //      64597 
       111: cosine = 18'b001111110001000100;  //      64580 
       112: cosine = 18'b001111110000110011;  //      64563 
       113: cosine = 18'b001111110000100001;  //      64545 
       114: cosine = 18'b001111110000010000;  //      64528 
       115: cosine = 18'b001111101111111110;  //      64510 
       116: cosine = 18'b001111101111101100;  //      64492 
       117: cosine = 18'b001111101111011010;  //      64474 
       118: cosine = 18'b001111101111001000;  //      64456 
       119: cosine = 18'b001111101110110110;  //      64438 
       120: cosine = 18'b001111101110100100;  //      64420 
       121: cosine = 18'b001111101110010001;  //      64401 
       122: cosine = 18'b001111101101111110;  //      64382 
       123: cosine = 18'b001111101101101011;  //      64363 
       124: cosine = 18'b001111101101011000;  //      64344 
       125: cosine = 18'b001111101101000101;  //      64325 
       126: cosine = 18'b001111101100110010;  //      64306 
       127: cosine = 18'b001111101100011111;  //      64287 
       128: cosine = 18'b001111101100001011;  //      64267 
       129: cosine = 18'b001111101011110111;  //      64247 
       130: cosine = 18'b001111101011100011;  //      64227 
       131: cosine = 18'b001111101011001111;  //      64207 
       132: cosine = 18'b001111101010111011;  //      64187 
       133: cosine = 18'b001111101010100111;  //      64167 
       134: cosine = 18'b001111101010010010;  //      64146 
       135: cosine = 18'b001111101001111101;  //      64125 
       136: cosine = 18'b001111101001101001;  //      64105 
       137: cosine = 18'b001111101001010100;  //      64084 
       138: cosine = 18'b001111101000111110;  //      64062 
       139: cosine = 18'b001111101000101001;  //      64041 
       140: cosine = 18'b001111101000010100;  //      64020 
       141: cosine = 18'b001111100111111110;  //      63998 
       142: cosine = 18'b001111100111101000;  //      63976 
       143: cosine = 18'b001111100111010011;  //      63955 
       144: cosine = 18'b001111100110111101;  //      63933 
       145: cosine = 18'b001111100110100110;  //      63910 
       146: cosine = 18'b001111100110010000;  //      63888 
       147: cosine = 18'b001111100101111010;  //      63866 
       148: cosine = 18'b001111100101100011;  //      63843 
       149: cosine = 18'b001111100101001100;  //      63820 
       150: cosine = 18'b001111100100110101;  //      63797 
       151: cosine = 18'b001111100100011110;  //      63774 
       152: cosine = 18'b001111100100000111;  //      63751 
       153: cosine = 18'b001111100011110000;  //      63728 
       154: cosine = 18'b001111100011011000;  //      63704 
       155: cosine = 18'b001111100011000000;  //      63680 
       156: cosine = 18'b001111100010101001;  //      63657 
       157: cosine = 18'b001111100010010001;  //      63633 
       158: cosine = 18'b001111100001111000;  //      63608 
       159: cosine = 18'b001111100001100000;  //      63584 
       160: cosine = 18'b001111100001001000;  //      63560 
       161: cosine = 18'b001111100000101111;  //      63535 
       162: cosine = 18'b001111100000010110;  //      63510 
       163: cosine = 18'b001111011111111110;  //      63486 
       164: cosine = 18'b001111011111100101;  //      63461 
       165: cosine = 18'b001111011111001011;  //      63435 
       166: cosine = 18'b001111011110110010;  //      63410 
       167: cosine = 18'b001111011110011001;  //      63385 
       168: cosine = 18'b001111011101111111;  //      63359 
       169: cosine = 18'b001111011101100101;  //      63333 
       170: cosine = 18'b001111011101001011;  //      63307 
       171: cosine = 18'b001111011100110001;  //      63281 
       172: cosine = 18'b001111011100010111;  //      63255 
       173: cosine = 18'b001111011011111101;  //      63229 
       174: cosine = 18'b001111011011100010;  //      63202 
       175: cosine = 18'b001111011011000111;  //      63175 
       176: cosine = 18'b001111011010101101;  //      63149 
       177: cosine = 18'b001111011010010010;  //      63122 
       178: cosine = 18'b001111011001110111;  //      63095 
       179: cosine = 18'b001111011001011011;  //      63067 
       180: cosine = 18'b001111011001000000;  //      63040 
       181: cosine = 18'b001111011000100100;  //      63012 
       182: cosine = 18'b001111011000001001;  //      62985 
       183: cosine = 18'b001111010111101101;  //      62957 
       184: cosine = 18'b001111010111010001;  //      62929 
       185: cosine = 18'b001111010110110101;  //      62901 
       186: cosine = 18'b001111010110011000;  //      62872 
       187: cosine = 18'b001111010101111100;  //      62844 
       188: cosine = 18'b001111010101011111;  //      62815 
       189: cosine = 18'b001111010101000011;  //      62787 
       190: cosine = 18'b001111010100100110;  //      62758 
       191: cosine = 18'b001111010100001001;  //      62729 
       192: cosine = 18'b001111010011101011;  //      62699 
       193: cosine = 18'b001111010011001110;  //      62670 
       194: cosine = 18'b001111010010110001;  //      62641 
       195: cosine = 18'b001111010010010011;  //      62611 
       196: cosine = 18'b001111010001110101;  //      62581 
       197: cosine = 18'b001111010001010111;  //      62551 
       198: cosine = 18'b001111010000111001;  //      62521 
       199: cosine = 18'b001111010000011011;  //      62491 
       200: cosine = 18'b001111001111111101;  //      62461 
       201: cosine = 18'b001111001111011110;  //      62430 
       202: cosine = 18'b001111001111000000;  //      62400 
       203: cosine = 18'b001111001110100001;  //      62369 
       204: cosine = 18'b001111001110000010;  //      62338 
       205: cosine = 18'b001111001101100011;  //      62307 
       206: cosine = 18'b001111001101000011;  //      62275 
       207: cosine = 18'b001111001100100100;  //      62244 
       208: cosine = 18'b001111001100000100;  //      62212 
       209: cosine = 18'b001111001011100101;  //      62181 
       210: cosine = 18'b001111001011000101;  //      62149 
       211: cosine = 18'b001111001010100101;  //      62117 
       212: cosine = 18'b001111001010000101;  //      62085 
       213: cosine = 18'b001111001001100101;  //      62053 
       214: cosine = 18'b001111001001000100;  //      62020 
       215: cosine = 18'b001111001000100100;  //      61988 
       216: cosine = 18'b001111001000000011;  //      61955 
       217: cosine = 18'b001111000111100010;  //      61922 
       218: cosine = 18'b001111000111000001;  //      61889 
       219: cosine = 18'b001111000110100000;  //      61856 
       220: cosine = 18'b001111000101111111;  //      61823 
       221: cosine = 18'b001111000101011101;  //      61789 
       222: cosine = 18'b001111000100111100;  //      61756 
       223: cosine = 18'b001111000100011010;  //      61722 
       224: cosine = 18'b001111000011111000;  //      61688 
       225: cosine = 18'b001111000011010110;  //      61654 
       226: cosine = 18'b001111000010110100;  //      61620 
       227: cosine = 18'b001111000010010010;  //      61586 
       228: cosine = 18'b001111000001101111;  //      61551 
       229: cosine = 18'b001111000001001101;  //      61517 
       230: cosine = 18'b001111000000101010;  //      61482 
       231: cosine = 18'b001111000000000111;  //      61447 
       232: cosine = 18'b001110111111100100;  //      61412 
       233: cosine = 18'b001110111111000001;  //      61377 
       234: cosine = 18'b001110111110011101;  //      61341 
       235: cosine = 18'b001110111101111010;  //      61306 
       236: cosine = 18'b001110111101010110;  //      61270 
       237: cosine = 18'b001110111100110011;  //      61235 
       238: cosine = 18'b001110111100001111;  //      61199 
       239: cosine = 18'b001110111011101011;  //      61163 
       240: cosine = 18'b001110111011000111;  //      61127 
       241: cosine = 18'b001110111010100010;  //      61090 
       242: cosine = 18'b001110111001111110;  //      61054 
       243: cosine = 18'b001110111001011001;  //      61017 
       244: cosine = 18'b001110111000110100;  //      60980 
       245: cosine = 18'b001110111000001111;  //      60943 
       246: cosine = 18'b001110110111101010;  //      60906 
       247: cosine = 18'b001110110111000101;  //      60869 
       248: cosine = 18'b001110110110100000;  //      60832 
       249: cosine = 18'b001110110101111010;  //      60794 
       250: cosine = 18'b001110110101010101;  //      60757 
       251: cosine = 18'b001110110100101111;  //      60719 
       252: cosine = 18'b001110110100001001;  //      60681 
       253: cosine = 18'b001110110011100011;  //      60643 
       254: cosine = 18'b001110110010111101;  //      60605 
       255: cosine = 18'b001110110010010111;  //      60567 
       256: cosine = 18'b001110110001110000;  //      60528 
       257: cosine = 18'b001110110001001010;  //      60490 
       258: cosine = 18'b001110110000100011;  //      60451 
       259: cosine = 18'b001110101111111100;  //      60412 
       260: cosine = 18'b001110101111010101;  //      60373 
       261: cosine = 18'b001110101110101110;  //      60334 
       262: cosine = 18'b001110101110000110;  //      60294 
       263: cosine = 18'b001110101101011111;  //      60255 
       264: cosine = 18'b001110101100110111;  //      60215 
       265: cosine = 18'b001110101100001111;  //      60175 
       266: cosine = 18'b001110101011101000;  //      60136 
       267: cosine = 18'b001110101011000000;  //      60096 
       268: cosine = 18'b001110101010010111;  //      60055 
       269: cosine = 18'b001110101001101111;  //      60015 
       270: cosine = 18'b001110101001000111;  //      59975 
       271: cosine = 18'b001110101000011110;  //      59934 
       272: cosine = 18'b001110100111110101;  //      59893 
       273: cosine = 18'b001110100111001100;  //      59852 
       274: cosine = 18'b001110100110100011;  //      59811 
       275: cosine = 18'b001110100101111010;  //      59770 
       276: cosine = 18'b001110100101010001;  //      59729 
       277: cosine = 18'b001110100100100111;  //      59687 
       278: cosine = 18'b001110100011111110;  //      59646 
       279: cosine = 18'b001110100011010100;  //      59604 
       280: cosine = 18'b001110100010101010;  //      59562 
       281: cosine = 18'b001110100010000000;  //      59520 
       282: cosine = 18'b001110100001010110;  //      59478 
       283: cosine = 18'b001110100000101100;  //      59436 
       284: cosine = 18'b001110100000000001;  //      59393 
       285: cosine = 18'b001110011111010111;  //      59351 
       286: cosine = 18'b001110011110101100;  //      59308 
       287: cosine = 18'b001110011110000001;  //      59265 
       288: cosine = 18'b001110011101010110;  //      59222 
       289: cosine = 18'b001110011100101011;  //      59179 
       290: cosine = 18'b001110011100000000;  //      59136 
       291: cosine = 18'b001110011011010101;  //      59093 
       292: cosine = 18'b001110011010101001;  //      59049 
       293: cosine = 18'b001110011001111101;  //      59005 
       294: cosine = 18'b001110011001010010;  //      58962 
       295: cosine = 18'b001110011000100110;  //      58918 
       296: cosine = 18'b001110010111111001;  //      58873 
       297: cosine = 18'b001110010111001101;  //      58829 
       298: cosine = 18'b001110010110100001;  //      58785 
       299: cosine = 18'b001110010101110100;  //      58740 
       300: cosine = 18'b001110010101001000;  //      58696 
       301: cosine = 18'b001110010100011011;  //      58651 
       302: cosine = 18'b001110010011101110;  //      58606 
       303: cosine = 18'b001110010011000001;  //      58561 
       304: cosine = 18'b001110010010010100;  //      58516 
       305: cosine = 18'b001110010001100110;  //      58470 
       306: cosine = 18'b001110010000111001;  //      58425 
       307: cosine = 18'b001110010000001011;  //      58379 
       308: cosine = 18'b001110001111011110;  //      58334 
       309: cosine = 18'b001110001110110000;  //      58288 
       310: cosine = 18'b001110001110000010;  //      58242 
       311: cosine = 18'b001110001101010011;  //      58195 
       312: cosine = 18'b001110001100100101;  //      58149 
       313: cosine = 18'b001110001011110111;  //      58103 
       314: cosine = 18'b001110001011001000;  //      58056 
       315: cosine = 18'b001110001010011001;  //      58009 
       316: cosine = 18'b001110001001101011;  //      57963 
       317: cosine = 18'b001110001000111100;  //      57916 
       318: cosine = 18'b001110001000001101;  //      57869 
       319: cosine = 18'b001110000111011101;  //      57821 
       320: cosine = 18'b001110000110101110;  //      57774 
       321: cosine = 18'b001110000101111110;  //      57726 
       322: cosine = 18'b001110000101001111;  //      57679 
       323: cosine = 18'b001110000100011111;  //      57631 
       324: cosine = 18'b001110000011101111;  //      57583 
       325: cosine = 18'b001110000010111111;  //      57535 
       326: cosine = 18'b001110000010001111;  //      57487 
       327: cosine = 18'b001110000001011110;  //      57438 
       328: cosine = 18'b001110000000101110;  //      57390 
       329: cosine = 18'b001101111111111101;  //      57341 
       330: cosine = 18'b001101111111001101;  //      57293 
       331: cosine = 18'b001101111110011100;  //      57244 
       332: cosine = 18'b001101111101101011;  //      57195 
       333: cosine = 18'b001101111100111001;  //      57145 
       334: cosine = 18'b001101111100001000;  //      57096 
       335: cosine = 18'b001101111011010111;  //      57047 
       336: cosine = 18'b001101111010100101;  //      56997 
       337: cosine = 18'b001101111001110100;  //      56948 
       338: cosine = 18'b001101111001000010;  //      56898 
       339: cosine = 18'b001101111000010000;  //      56848 
       340: cosine = 18'b001101110111011110;  //      56798 
       341: cosine = 18'b001101110110101011;  //      56747 
       342: cosine = 18'b001101110101111001;  //      56697 
       343: cosine = 18'b001101110101000111;  //      56647 
       344: cosine = 18'b001101110100010100;  //      56596 
       345: cosine = 18'b001101110011100001;  //      56545 
       346: cosine = 18'b001101110010101110;  //      56494 
       347: cosine = 18'b001101110001111011;  //      56443 
       348: cosine = 18'b001101110001001000;  //      56392 
       349: cosine = 18'b001101110000010101;  //      56341 
       350: cosine = 18'b001101101111100001;  //      56289 
       351: cosine = 18'b001101101110101110;  //      56238 
       352: cosine = 18'b001101101101111010;  //      56186 
       353: cosine = 18'b001101101101000110;  //      56134 
       354: cosine = 18'b001101101100010010;  //      56082 
       355: cosine = 18'b001101101011011110;  //      56030 
       356: cosine = 18'b001101101010101010;  //      55978 
       357: cosine = 18'b001101101001110110;  //      55926 
       358: cosine = 18'b001101101001000001;  //      55873 
       359: cosine = 18'b001101101000001101;  //      55821 
       360: cosine = 18'b001101100111011000;  //      55768 
       361: cosine = 18'b001101100110100011;  //      55715 
       362: cosine = 18'b001101100101101110;  //      55662 
       363: cosine = 18'b001101100100111001;  //      55609 
       364: cosine = 18'b001101100100000100;  //      55556 
       365: cosine = 18'b001101100011001110;  //      55502 
       366: cosine = 18'b001101100010011001;  //      55449 
       367: cosine = 18'b001101100001100011;  //      55395 
       368: cosine = 18'b001101100000101101;  //      55341 
       369: cosine = 18'b001101011111111000;  //      55288 
       370: cosine = 18'b001101011111000001;  //      55233 
       371: cosine = 18'b001101011110001011;  //      55179 
       372: cosine = 18'b001101011101010101;  //      55125 
       373: cosine = 18'b001101011100011111;  //      55071 
       374: cosine = 18'b001101011011101000;  //      55016 
       375: cosine = 18'b001101011010110001;  //      54961 
       376: cosine = 18'b001101011001111010;  //      54906 
       377: cosine = 18'b001101011001000100;  //      54852 
       378: cosine = 18'b001101011000001100;  //      54796 
       379: cosine = 18'b001101010111010101;  //      54741 
       380: cosine = 18'b001101010110011110;  //      54686 
       381: cosine = 18'b001101010101100110;  //      54630 
       382: cosine = 18'b001101010100101111;  //      54575 
       383: cosine = 18'b001101010011110111;  //      54519 
       384: cosine = 18'b001101010010111111;  //      54463 
       385: cosine = 18'b001101010010000111;  //      54407 
       386: cosine = 18'b001101010001001111;  //      54351 
       387: cosine = 18'b001101010000010111;  //      54295 
       388: cosine = 18'b001101001111011111;  //      54239 
       389: cosine = 18'b001101001110100110;  //      54182 
       390: cosine = 18'b001101001101101101;  //      54125 
       391: cosine = 18'b001101001100110101;  //      54069 
       392: cosine = 18'b001101001011111100;  //      54012 
       393: cosine = 18'b001101001011000011;  //      53955 
       394: cosine = 18'b001101001010001010;  //      53898 
       395: cosine = 18'b001101001001010000;  //      53840 
       396: cosine = 18'b001101001000010111;  //      53783 
       397: cosine = 18'b001101000111011110;  //      53726 
       398: cosine = 18'b001101000110100100;  //      53668 
       399: cosine = 18'b001101000101101010;  //      53610 
       400: cosine = 18'b001101000100110000;  //      53552 
       401: cosine = 18'b001101000011110110;  //      53494 
       402: cosine = 18'b001101000010111100;  //      53436 
       403: cosine = 18'b001101000010000010;  //      53378 
       404: cosine = 18'b001101000001000111;  //      53319 
       405: cosine = 18'b001101000000001101;  //      53261 
       406: cosine = 18'b001100111111010010;  //      53202 
       407: cosine = 18'b001100111110011000;  //      53144 
       408: cosine = 18'b001100111101011101;  //      53085 
       409: cosine = 18'b001100111100100010;  //      53026 
       410: cosine = 18'b001100111011100111;  //      52967 
       411: cosine = 18'b001100111010101011;  //      52907 
       412: cosine = 18'b001100111001110000;  //      52848 
       413: cosine = 18'b001100111000110100;  //      52788 
       414: cosine = 18'b001100110111111001;  //      52729 
       415: cosine = 18'b001100110110111101;  //      52669 
       416: cosine = 18'b001100110110000001;  //      52609 
       417: cosine = 18'b001100110101000101;  //      52549 
       418: cosine = 18'b001100110100001001;  //      52489 
       419: cosine = 18'b001100110011001101;  //      52429 
       420: cosine = 18'b001100110010010000;  //      52368 
       421: cosine = 18'b001100110001010100;  //      52308 
       422: cosine = 18'b001100110000010111;  //      52247 
       423: cosine = 18'b001100101111011010;  //      52186 
       424: cosine = 18'b001100101110011110;  //      52126 
       425: cosine = 18'b001100101101100001;  //      52065 
       426: cosine = 18'b001100101100100011;  //      52003 
       427: cosine = 18'b001100101011100110;  //      51942 
       428: cosine = 18'b001100101010101001;  //      51881 
       429: cosine = 18'b001100101001101011;  //      51819 
       430: cosine = 18'b001100101000101110;  //      51758 
       431: cosine = 18'b001100100111110000;  //      51696 
       432: cosine = 18'b001100100110110010;  //      51634 
       433: cosine = 18'b001100100101110100;  //      51572 
       434: cosine = 18'b001100100100110110;  //      51510 
       435: cosine = 18'b001100100011111000;  //      51448 
       436: cosine = 18'b001100100010111010;  //      51386 
       437: cosine = 18'b001100100001111011;  //      51323 
       438: cosine = 18'b001100100000111100;  //      51260 
       439: cosine = 18'b001100011111111110;  //      51198 
       440: cosine = 18'b001100011110111111;  //      51135 
       441: cosine = 18'b001100011110000000;  //      51072 
       442: cosine = 18'b001100011101000001;  //      51009 
       443: cosine = 18'b001100011100000010;  //      50946 
       444: cosine = 18'b001100011011000010;  //      50882 
       445: cosine = 18'b001100011010000011;  //      50819 
       446: cosine = 18'b001100011001000100;  //      50756 
       447: cosine = 18'b001100011000000100;  //      50692 
       448: cosine = 18'b001100010111000100;  //      50628 
       449: cosine = 18'b001100010110000100;  //      50564 
       450: cosine = 18'b001100010101000100;  //      50500 
       451: cosine = 18'b001100010100000100;  //      50436 
       452: cosine = 18'b001100010011000100;  //      50372 
       453: cosine = 18'b001100010010000011;  //      50307 
       454: cosine = 18'b001100010001000011;  //      50243 
       455: cosine = 18'b001100010000000010;  //      50178 
       456: cosine = 18'b001100001111000010;  //      50114 
       457: cosine = 18'b001100001110000001;  //      50049 
       458: cosine = 18'b001100001101000000;  //      49984 
       459: cosine = 18'b001100001011111111;  //      49919 
       460: cosine = 18'b001100001010111110;  //      49854 
       461: cosine = 18'b001100001001111100;  //      49788 
       462: cosine = 18'b001100001000111011;  //      49723 
       463: cosine = 18'b001100000111111001;  //      49657 
       464: cosine = 18'b001100000110111000;  //      49592 
       465: cosine = 18'b001100000101110110;  //      49526 
       466: cosine = 18'b001100000100110100;  //      49460 
       467: cosine = 18'b001100000011110010;  //      49394 
       468: cosine = 18'b001100000010110000;  //      49328 
       469: cosine = 18'b001100000001101110;  //      49262 
       470: cosine = 18'b001100000000101011;  //      49195 
       471: cosine = 18'b001011111111101001;  //      49129 
       472: cosine = 18'b001011111110100110;  //      49062 
       473: cosine = 18'b001011111101100011;  //      48995 
       474: cosine = 18'b001011111100100001;  //      48929 
       475: cosine = 18'b001011111011011110;  //      48862 
       476: cosine = 18'b001011111010011011;  //      48795 
       477: cosine = 18'b001011111001010111;  //      48727 
       478: cosine = 18'b001011111000010100;  //      48660 
       479: cosine = 18'b001011110111010001;  //      48593 
       480: cosine = 18'b001011110110001101;  //      48525 
       481: cosine = 18'b001011110101001010;  //      48458 
       482: cosine = 18'b001011110100000110;  //      48390 
       483: cosine = 18'b001011110011000010;  //      48322 
       484: cosine = 18'b001011110001111110;  //      48254 
       485: cosine = 18'b001011110000111010;  //      48186 
       486: cosine = 18'b001011101111110110;  //      48118 
       487: cosine = 18'b001011101110110001;  //      48049 
       488: cosine = 18'b001011101101101101;  //      47981 
       489: cosine = 18'b001011101100101000;  //      47912 
       490: cosine = 18'b001011101011100100;  //      47844 
       491: cosine = 18'b001011101010011111;  //      47775 
       492: cosine = 18'b001011101001011010;  //      47706 
       493: cosine = 18'b001011101000010101;  //      47637 
       494: cosine = 18'b001011100111010000;  //      47568 
       495: cosine = 18'b001011100110001011;  //      47499 
       496: cosine = 18'b001011100101000110;  //      47430 
       497: cosine = 18'b001011100100000000;  //      47360 
       498: cosine = 18'b001011100010111011;  //      47291 
       499: cosine = 18'b001011100001110101;  //      47221 
       500: cosine = 18'b001011100000101111;  //      47151 
       501: cosine = 18'b001011011111101001;  //      47081 
       502: cosine = 18'b001011011110100011;  //      47011 
       503: cosine = 18'b001011011101011101;  //      46941 
       504: cosine = 18'b001011011100010111;  //      46871 
       505: cosine = 18'b001011011011010001;  //      46801 
       506: cosine = 18'b001011011010001010;  //      46730 
       507: cosine = 18'b001011011001000100;  //      46660 
       508: cosine = 18'b001011010111111101;  //      46589 
       509: cosine = 18'b001011010110110110;  //      46518 
       510: cosine = 18'b001011010101101111;  //      46447 
       511: cosine = 18'b001011010100101000;  //      46376 
    endcase 
endmodule 


