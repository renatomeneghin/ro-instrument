`timescale 1ns/10ps

module COREFFT_C0_COREFFT_C0_0_twidLut_stage_2 (index, twid_im, twid_re);
  input[9:0] index;
  output [31:0] twid_im, twid_re;
  reg    signed [31:0] twid_im, twid_re;

  always @ (index) 
    case (index) 
   0 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   1 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   2 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   3 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   4 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   5 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   6 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   7 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   8 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   9 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  10 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  11 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  12 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  13 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  14 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  15 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  16 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  17 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  18 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  19 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  20 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  21 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  22 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  23 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  24 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  25 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  26 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  27 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  28 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  29 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  30 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  31 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  32 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  33 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  34 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  35 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  36 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  37 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  38 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  39 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  40 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  41 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  42 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  43 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  44 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  45 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  46 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  47 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  48 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  49 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  50 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  51 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  52 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  53 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  54 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  55 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  56 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  57 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  58 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  59 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  60 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  61 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  62 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  63 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  64 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  65 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  66 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  67 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  68 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  69 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  70 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  71 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  72 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  73 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  74 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  75 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  76 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  77 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  78 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  79 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  80 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  81 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  82 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  83 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  84 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  85 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  86 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  87 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  88 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  89 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  90 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  91 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  92 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  93 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  94 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  95 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  96 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  97 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  98 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  99 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 100 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 101 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 102 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 103 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 104 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 105 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 106 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 107 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 108 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 109 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 110 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 111 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 112 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 113 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 114 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 115 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 116 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 117 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 118 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 119 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 120 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 121 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 122 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 123 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 124 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 125 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 126 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 127 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 128 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 129 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 130 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 131 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 132 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 133 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 134 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 135 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 136 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 137 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 138 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 139 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 140 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 141 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 142 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 143 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 144 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 145 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 146 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 147 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 148 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 149 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 150 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 151 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 152 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 153 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 154 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 155 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 156 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 157 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 158 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 159 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 160 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 161 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 162 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 163 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 164 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 165 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 166 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 167 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 168 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 169 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 170 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 171 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 172 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 173 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 174 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 175 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 176 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 177 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 178 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 179 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 180 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 181 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 182 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 183 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 184 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 185 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 186 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 187 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 188 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 189 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 190 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 191 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 192 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 193 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 194 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 195 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 196 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 197 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 198 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 199 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 200 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 201 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 202 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 203 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 204 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 205 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 206 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 207 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 208 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 209 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 210 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 211 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 212 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 213 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 214 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 215 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 216 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 217 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 218 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 219 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 220 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 221 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 222 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 223 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 224 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 225 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 226 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 227 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 228 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 229 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 230 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 231 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 232 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 233 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 234 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 235 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 236 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 237 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 238 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 239 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 240 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 241 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 242 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 243 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 244 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 245 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 246 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 247 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 248 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 249 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 250 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 251 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 252 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 253 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 254 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 255 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 256 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 257 : begin twid_im = 32'b11111110011011011110001011100000; twid_re = 32'b01111111111111011000100001011001; end  //-0,012  1,000
 258 : begin twid_im = 32'b11111100110110111101010101000001; twid_re = 32'b01111111111101100010000110000001; end  //-0,025  1,000
 259 : begin twid_im = 32'b11111011010010011110011010100011; twid_re = 32'b01111111111010011100101110111111; end  //-0,037  0,999
 260 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b01111111110110001000011110001101; end  //-0,049  0,999
 261 : begin twid_im = 32'b11111000001001101010010001100010; twid_re = 32'b01111111110000100101010110010101; end  //-0,061  0,998
 262 : begin twid_im = 32'b11110110100101010110111110110111; twid_re = 32'b01111111101001110011011010110011; end  //-0,074  0,997
 263 : begin twid_im = 32'b11110101000001001001011111111011; twid_re = 32'b01111111100001110010101111110010; end  //-0,086  0,996
 264 : begin twid_im = 32'b11110011011101000010110010100010; twid_re = 32'b01111111011000100011011010001110; end  //-0,098  0,995
 265 : begin twid_im = 32'b11110001111001000011110100011100; twid_re = 32'b01111111001110000101011111110101; end  //-0,110  0,994
 266 : begin twid_im = 32'b11110000010101001101100011010101; twid_re = 32'b01111111000010011001000111000011; end  //-0,122  0,992
 267 : begin twid_im = 32'b11101110110001100000111100110001; twid_re = 32'b01111110110101011110010111000101; end  //-0,135  0,991
 268 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b01111110100111010101010111111011; end  //-0,147  0,989
 269 : begin twid_im = 32'b11101011101010101000100101001111; twid_re = 32'b01111110010111111110010010010010; end  //-0,159  0,987
 270 : begin twid_im = 32'b11101010000111011110101110111100; twid_re = 32'b01111110000111011001001111101001; end  //-0,171  0,985
 271 : begin twid_im = 32'b11101000100100100010011000100010; twid_re = 32'b01111101110101100110011010001110; end  //-0,183  0,983
 272 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b01111101100010100101111100111111; end  //-0,195  0,981
 273 : begin twid_im = 32'b11100101011111010101111111011011; twid_re = 32'b01111101001110011000000011101011; end  //-0,207  0,978
 274 : begin twid_im = 32'b11100011111101000111110110010110; twid_re = 32'b01111100111000111100111010110001; end  //-0,219  0,976
 275 : begin twid_im = 32'b11100010011011001011000000011011; twid_re = 32'b01111100100010010100101111011101; end  //-0,231  0,973
 276 : begin twid_im = 32'b11100000111001100000011010000101; twid_re = 32'b01111100001010011111101111101101; end  //-0,243  0,970
 277 : begin twid_im = 32'b11011111011000001000111111100100; twid_re = 32'b01111011110001011110001010001111; end  //-0,255  0,967
 278 : begin twid_im = 32'b11011101110111000101101100111011; twid_re = 32'b01111011010111010000001110011101; end  //-0,267  0,964
 279 : begin twid_im = 32'b11011100010110010111011110000010; twid_re = 32'b01111010111011110110001100100011; end  //-0,279  0,960
 280 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
 281 : begin twid_im = 32'b11011001010101111101111001111011; twid_re = 32'b01111010000001011110111010101100; end  //-0,302  0,953
 282 : begin twid_im = 32'b11010111110110010100011011011000; twid_re = 32'b01111001100010100010001110110000; end  //-0,314  0,950
 283 : begin twid_im = 32'b11010110010111000011101101111011; twid_re = 32'b01111001000010011010100100101100; end  //-0,325  0,946
 284 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b01111000100001001000010000010011; end  //-0,337  0,942
 285 : begin twid_im = 32'b11010011011001110000010001000110; twid_re = 32'b01110111111110101011100110001000; end  //-0,348  0,937
 286 : begin twid_im = 32'b11010001111011101111010110011110; twid_re = 32'b01110111011011000100111011011010; end  //-0,360  0,933
 287 : begin twid_im = 32'b11010000011110001010110110011110; twid_re = 32'b01110110110110010100100110001000; end  //-0,371  0,929
 288 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b01110110010000011010111100111100; end  //-0,383  0,924
 289 : begin twid_im = 32'b11001101100100011010101100111001; twid_re = 32'b01110101101001011000010111001110; end  //-0,394  0,919
 290 : begin twid_im = 32'b11001100001000010000110101111001; twid_re = 32'b01110101000001001101001101000100; end  //-0,405  0,914
 291 : begin twid_im = 32'b11001010101100100110111110101010; twid_re = 32'b01110100010111111001110111010000; end  //-0,416  0,909
 292 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b01110011101101011110101111010000; end  //-0,428  0,904
 293 : begin twid_im = 32'b11000111110110110110110001010000; twid_re = 32'b01110011000001111100001111001111; end  //-0,439  0,899
 294 : begin twid_im = 32'b11000110011100110010001011001110; twid_re = 32'b01110010010101010010110010000100; end  //-0,450  0,893
 295 : begin twid_im = 32'b11000101000011010001000101001001; twid_re = 32'b01110001100111100010110011010001; end  //-0,461  0,888
 296 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b01110000111000101100101111000101; end  //-0,471  0,882
 297 : begin twid_im = 32'b11000010010001111100110101011011; twid_re = 32'b01110000001000110001000010011001; end  //-0,482  0,876
 298 : begin twid_im = 32'b11000000111010001011011001001001; twid_re = 32'b01101111010111110000001010110001; end  //-0,493  0,870
 299 : begin twid_im = 32'b10111111100011000000110111100011; twid_re = 32'b01101110100101101010100110011100; end  //-0,504  0,864
 300 : begin twid_im = 32'b10111110001100011110000110011100; twid_re = 32'b01101101110010100000110100010100; end  //-0,514  0,858
 301 : begin twid_im = 32'b10111100110110100011111011001011; twid_re = 32'b01101100111110010011010011111011; end  //-0,525  0,851
 302 : begin twid_im = 32'b10111011100001010011001010110000; twid_re = 32'b01101100001001000010100101011111; end  //-0,535  0,845
 303 : begin twid_im = 32'b10111010001100101100101001110001; twid_re = 32'b01101011010010101111001001111000; end  //-0,545  0,838
 304 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
 305 : begin twid_im = 32'b10110111100101100001100110011100; twid_re = 32'b01101001100011000010010001101011; end  //-0,566  0,825
 306 : begin twid_im = 32'b10110110010010111110101011001101; twid_re = 32'b01101000101001101001111010000000; end  //-0,576  0,818
 307 : begin twid_im = 32'b10110101000001001001001101101001; twid_re = 32'b01100111101111010000111110111100; end  //-0,586  0,810
 308 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b01100110110011111000000100011111; end  //-0,596  0,803
 309 : begin twid_im = 32'b10110010011111101001110100111101; twid_re = 32'b01100101110111011111101111010010; end  //-0,606  0,796
 310 : begin twid_im = 32'b10110001010000000001011101011100; twid_re = 32'b01100100111010001000100100100101; end  //-0,615  0,788
 311 : begin twid_im = 32'b10110000000001001001101010110100; twid_re = 32'b01100011111011110011001010001111; end  //-0,625  0,781
 312 : begin twid_im = 32'b10101110110011000011001101101100; twid_re = 32'b01100010111100100000000110101100; end  //-0,634  0,773
 313 : begin twid_im = 32'b10101101100101101110110110010010; twid_re = 32'b01100001111100010000000000111110; end  //-0,644  0,765
 314 : begin twid_im = 32'b10101100011001001101010100010001; twid_re = 32'b01100000111011000011100000101111; end  //-0,653  0,757
 315 : begin twid_im = 32'b10101011001101011111010110110110; twid_re = 32'b01011111111000111011001110001101; end  //-0,662  0,749
 316 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b01011110110101110111110010001001; end  //-0,672  0,741
 317 : begin twid_im = 32'b10101000111000100001000100000111; twid_re = 32'b01011101110001111001110101111011; end  //-0,681  0,733
 318 : begin twid_im = 32'b10100111101111010010001010101100; twid_re = 32'b01011100101101000010000011011111; end  //-0,690  0,724
 319 : begin twid_im = 32'b10100110100110111001101101101001; twid_re = 32'b01011011100111010001000101010011; end  //-0,698  0,716
 320 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
 321 : begin twid_im = 32'b10100100011000101110111010101101; twid_re = 32'b01011001011001000110010010010111; end  //-0,716  0,698
 322 : begin twid_im = 32'b10100011010010111101111100100001; twid_re = 32'b01011000010000101101110101010100; end  //-0,724  0,690
 323 : begin twid_im = 32'b10100010001110000110001010000101; twid_re = 32'b01010111000111011110111011111001; end  //-0,733  0,681
 324 : begin twid_im = 32'b10100001001010001000001101110111; twid_re = 32'b01010101111101011010010011010010; end  //-0,741  0,672
 325 : begin twid_im = 32'b10100000000111000100110001110011; twid_re = 32'b01010100110010100000101001001010; end  //-0,749  0,662
 326 : begin twid_im = 32'b10011111000100111100011111010001; twid_re = 32'b01010011100110110010101011101111; end  //-0,757  0,653
 327 : begin twid_im = 32'b10011110000011101111111111000010; twid_re = 32'b01010010011010010001001001101110; end  //-0,765  0,644
 328 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
 329 : begin twid_im = 32'b10011100000100001100110101110001; twid_re = 32'b01001111111110110110010101001100; end  //-0,781  0,625
 330 : begin twid_im = 32'b10011011000101110111011011011011; twid_re = 32'b01001110101111111110100010100100; end  //-0,788  0,615
 331 : begin twid_im = 32'b10011010001000100000010000101110; twid_re = 32'b01001101100000010110001011000011; end  //-0,796  0,606
 332 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b01001100001111111101111111110011; end  //-0,803  0,596
 333 : begin twid_im = 32'b10011000010000101111000001000100; twid_re = 32'b01001010111110110110110010010111; end  //-0,810  0,586
 334 : begin twid_im = 32'b10010111010110010110000110000000; twid_re = 32'b01001001101101000001010100110011; end  //-0,818  0,576
 335 : begin twid_im = 32'b10010110011100111101101110010101; twid_re = 32'b01001000011010011110011001100100; end  //-0,825  0,566
 336 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b01000111000111001110110011100110; end  //-0,831  0,556
 337 : begin twid_im = 32'b10010100101101010000110110001000; twid_re = 32'b01000101110011010011010110001111; end  //-0,838  0,545
 338 : begin twid_im = 32'b10010011110110111101011010100001; twid_re = 32'b01000100011110101100110101010000; end  //-0,845  0,535
 339 : begin twid_im = 32'b10010011000001101100101100000101; twid_re = 32'b01000011001001011100000100110101; end  //-0,851  0,525
 340 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b01000001110011100001111001100100; end  //-0,858  0,514
 341 : begin twid_im = 32'b10010001011010010101011001100100; twid_re = 32'b01000000011100111111001000011101; end  //-0,864  0,504
 342 : begin twid_im = 32'b10010000101000001111110101001111; twid_re = 32'b00111111000101110100100110110111; end  //-0,870  0,493
 343 : begin twid_im = 32'b10001111110111001110111101100111; twid_re = 32'b00111101101110000011001010100101; end  //-0,876  0,482
 344 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b00111100010101101011101001110000; end  //-0,882  0,471
 345 : begin twid_im = 32'b10001110011000011101001100101111; twid_re = 32'b00111010111100101110111010110111; end  //-0,888  0,461
 346 : begin twid_im = 32'b10001101101010101101001101111100; twid_re = 32'b00111001100011001101110100110010; end  //-0,893  0,450
 347 : begin twid_im = 32'b10001100111110000011110000110001; twid_re = 32'b00111000001001001001001110110000; end  //-0,899  0,439
 348 : begin twid_im = 32'b10001100010010100001010000110000; twid_re = 32'b00110110101110100010000000010011; end  //-0,904  0,428
 349 : begin twid_im = 32'b10001011101000000110001000110000; twid_re = 32'b00110101010011011001000001010110; end  //-0,909  0,416
 350 : begin twid_im = 32'b10001010111110110010110010111100; twid_re = 32'b00110011110111101111001010000111; end  //-0,914  0,405
 351 : begin twid_im = 32'b10001010010110100111101000110010; twid_re = 32'b00110010011011100101010011000111; end  //-0,919  0,394
 352 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
 353 : begin twid_im = 32'b10001001001001101011011001111000; twid_re = 32'b00101111100001110101001001100010; end  //-0,929  0,371
 354 : begin twid_im = 32'b10001000100100111011000100100110; twid_re = 32'b00101110000100010000101001100010; end  //-0,933  0,360
 355 : begin twid_im = 32'b10001000000001010100011001111000; twid_re = 32'b00101100100110001111101110111010; end  //-0,937  0,348
 356 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b00101011000111110011010011101011; end  //-0,942  0,337
 357 : begin twid_im = 32'b10000110111101100101011011010100; twid_re = 32'b00101001101000111100010010000101; end  //-0,946  0,325
 358 : begin twid_im = 32'b10000110011101011101110001010000; twid_re = 32'b00101000001001101011100100101000; end  //-0,950  0,314
 359 : begin twid_im = 32'b10000101111110100001000101010100; twid_re = 32'b00100110101010000010000110000101; end  //-0,953  0,302
 360 : begin twid_im = 32'b10000101100000101111101010100110; twid_re = 32'b00100101001010000000110001011101; end  //-0,957  0,290
 361 : begin twid_im = 32'b10000101000100001001110011011101; twid_re = 32'b00100011101001101000100001111110; end  //-0,960  0,279
 362 : begin twid_im = 32'b10000100101000101111110001100011; twid_re = 32'b00100010001000111010010011000101; end  //-0,964  0,267
 363 : begin twid_im = 32'b10000100001110100001110101110001; twid_re = 32'b00100000100111110111000000011100; end  //-0,967  0,255
 364 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b00011111000110011111100101111011; end  //-0,970  0,243
 365 : begin twid_im = 32'b10000011011101101011010000100011; twid_re = 32'b00011101100100110100111111100101; end  //-0,973  0,231
 366 : begin twid_im = 32'b10000011000111000011000101001111; twid_re = 32'b00011100000010111000001001101010; end  //-0,976  0,219
 367 : begin twid_im = 32'b10000010110001100111111100010101; twid_re = 32'b00011010100000101010000000100101; end  //-0,978  0,207
 368 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b00011000111110001011100000111100; end  //-0,981  0,195
 369 : begin twid_im = 32'b10000010001010011001100101110010; twid_re = 32'b00010111011011011101100111011110; end  //-0,983  0,183
 370 : begin twid_im = 32'b10000001111000100110110000010111; twid_re = 32'b00010101111000100001010001000100; end  //-0,985  0,171
 371 : begin twid_im = 32'b10000001101000000001101101101110; twid_re = 32'b00010100010101010111011010110001; end  //-0,987  0,159
 372 : begin twid_im = 32'b10000001011000101010101000000101; twid_re = 32'b00010010110010000001000001101110; end  //-0,989  0,147
 373 : begin twid_im = 32'b10000001001010100001101000111011; twid_re = 32'b00010001001110011111000011001111; end  //-0,991  0,135
 374 : begin twid_im = 32'b10000000111101100110111000111101; twid_re = 32'b00001111101010110010011100101011; end  //-0,992  0,122
 375 : begin twid_im = 32'b10000000110001111010100000001011; twid_re = 32'b00001110000110111100001011100100; end  //-0,994  0,110
 376 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
 377 : begin twid_im = 32'b10000000011110001101010000001110; twid_re = 32'b00001010111110110110100000000101; end  //-0,996  0,086
 378 : begin twid_im = 32'b10000000010110001100100101001101; twid_re = 32'b00001001011010101001000001001001; end  //-0,997  0,074
 379 : begin twid_im = 32'b10000000001111011010101001101011; twid_re = 32'b00000111110110010101101110011110; end  //-0,998  0,061
 380 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b00000110010001111101100101111100; end  //-0,999  0,049
 381 : begin twid_im = 32'b10000000000101100011010001000001; twid_re = 32'b00000100101101100001100101011101; end  //-0,999  0,037
 382 : begin twid_im = 32'b10000000000010011101111001111111; twid_re = 32'b00000011001001000010101010111111; end  //-1,000  0,025
 383 : begin twid_im = 32'b10000000000000100111011110100111; twid_re = 32'b00000001100100100001110100100000; end  //-1,000  0,012
 384 : begin twid_im = 32'b10000000000000000000000000000001; twid_re = 32'b00000000000000000000000000000000; end  //-1,000  0,000
 385 : begin twid_im = 32'b10000000000000100111011110100111; twid_re = 32'b11111110011011011110001011100000; end  //-1,000 -0,012
 386 : begin twid_im = 32'b10000000000010011101111001111111; twid_re = 32'b11111100110110111101010101000001; end  //-1,000 -0,025
 387 : begin twid_im = 32'b10000000000101100011010001000001; twid_re = 32'b11111011010010011110011010100011; end  //-0,999 -0,037
 388 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b11111001101110000010011010000100; end  //-0,999 -0,049
 389 : begin twid_im = 32'b10000000001111011010101001101011; twid_re = 32'b11111000001001101010010001100010; end  //-0,998 -0,061
 390 : begin twid_im = 32'b10000000010110001100100101001101; twid_re = 32'b11110110100101010110111110110111; end  //-0,997 -0,074
 391 : begin twid_im = 32'b10000000011110001101010000001110; twid_re = 32'b11110101000001001001011111111011; end  //-0,996 -0,086
 392 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b11110011011101000010110010100010; end  //-0,995 -0,098
 393 : begin twid_im = 32'b10000000110001111010100000001011; twid_re = 32'b11110001111001000011110100011100; end  //-0,994 -0,110
 394 : begin twid_im = 32'b10000000111101100110111000111101; twid_re = 32'b11110000010101001101100011010101; end  //-0,992 -0,122
 395 : begin twid_im = 32'b10000001001010100001101000111011; twid_re = 32'b11101110110001100000111100110001; end  //-0,991 -0,135
 396 : begin twid_im = 32'b10000001011000101010101000000101; twid_re = 32'b11101101001101111110111110010010; end  //-0,989 -0,147
 397 : begin twid_im = 32'b10000001101000000001101101101110; twid_re = 32'b11101011101010101000100101001111; end  //-0,987 -0,159
 398 : begin twid_im = 32'b10000001111000100110110000010111; twid_re = 32'b11101010000111011110101110111100; end  //-0,985 -0,171
 399 : begin twid_im = 32'b10000010001010011001100101110010; twid_re = 32'b11101000100100100010011000100010; end  //-0,983 -0,183
 400 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b11100111000001110100011111000100; end  //-0,981 -0,195
 401 : begin twid_im = 32'b10000010110001100111111100010101; twid_re = 32'b11100101011111010101111111011011; end  //-0,978 -0,207
 402 : begin twid_im = 32'b10000011000111000011000101001111; twid_re = 32'b11100011111101000111110110010110; end  //-0,976 -0,219
 403 : begin twid_im = 32'b10000011011101101011010000100011; twid_re = 32'b11100010011011001011000000011011; end  //-0,973 -0,231
 404 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b11100000111001100000011010000101; end  //-0,970 -0,243
 405 : begin twid_im = 32'b10000100001110100001110101110001; twid_re = 32'b11011111011000001000111111100100; end  //-0,967 -0,255
 406 : begin twid_im = 32'b10000100101000101111110001100011; twid_re = 32'b11011101110111000101101100111011; end  //-0,964 -0,267
 407 : begin twid_im = 32'b10000101000100001001110011011101; twid_re = 32'b11011100010110010111011110000010; end  //-0,960 -0,279
 408 : begin twid_im = 32'b10000101100000101111101010100110; twid_re = 32'b11011010110101111111001110100011; end  //-0,957 -0,290
 409 : begin twid_im = 32'b10000101111110100001000101010100; twid_re = 32'b11011001010101111101111001111011; end  //-0,953 -0,302
 410 : begin twid_im = 32'b10000110011101011101110001010000; twid_re = 32'b11010111110110010100011011011000; end  //-0,950 -0,314
 411 : begin twid_im = 32'b10000110111101100101011011010100; twid_re = 32'b11010110010111000011101101111011; end  //-0,946 -0,325
 412 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b11010100111000001100101100010101; end  //-0,942 -0,337
 413 : begin twid_im = 32'b10001000000001010100011001111000; twid_re = 32'b11010011011001110000010001000110; end  //-0,937 -0,348
 414 : begin twid_im = 32'b10001000100100111011000100100110; twid_re = 32'b11010001111011101111010110011110; end  //-0,933 -0,360
 415 : begin twid_im = 32'b10001001001001101011011001111000; twid_re = 32'b11010000011110001010110110011110; end  //-0,929 -0,371
 416 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b11001111000001000011101010110011; end  //-0,924 -0,383
 417 : begin twid_im = 32'b10001010010110100111101000110010; twid_re = 32'b11001101100100011010101100111001; end  //-0,919 -0,394
 418 : begin twid_im = 32'b10001010111110110010110010111100; twid_re = 32'b11001100001000010000110101111001; end  //-0,914 -0,405
 419 : begin twid_im = 32'b10001011101000000110001000110000; twid_re = 32'b11001010101100100110111110101010; end  //-0,909 -0,416
 420 : begin twid_im = 32'b10001100010010100001010000110000; twid_re = 32'b11001001010001011101111111101101; end  //-0,904 -0,428
 421 : begin twid_im = 32'b10001100111110000011110000110001; twid_re = 32'b11000111110110110110110001010000; end  //-0,899 -0,439
 422 : begin twid_im = 32'b10001101101010101101001101111100; twid_re = 32'b11000110011100110010001011001110; end  //-0,893 -0,450
 423 : begin twid_im = 32'b10001110011000011101001100101111; twid_re = 32'b11000101000011010001000101001001; end  //-0,888 -0,461
 424 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b11000011101010010100010110010000; end  //-0,882 -0,471
 425 : begin twid_im = 32'b10001111110111001110111101100111; twid_re = 32'b11000010010001111100110101011011; end  //-0,876 -0,482
 426 : begin twid_im = 32'b10010000101000001111110101001111; twid_re = 32'b11000000111010001011011001001001; end  //-0,870 -0,493
 427 : begin twid_im = 32'b10010001011010010101011001100100; twid_re = 32'b10111111100011000000110111100011; end  //-0,864 -0,504
 428 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b10111110001100011110000110011100; end  //-0,858 -0,514
 429 : begin twid_im = 32'b10010011000001101100101100000101; twid_re = 32'b10111100110110100011111011001011; end  //-0,851 -0,525
 430 : begin twid_im = 32'b10010011110110111101011010100001; twid_re = 32'b10111011100001010011001010110000; end  //-0,845 -0,535
 431 : begin twid_im = 32'b10010100101101010000110110001000; twid_re = 32'b10111010001100101100101001110001; end  //-0,838 -0,545
 432 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b10111000111000110001001100011010; end  //-0,831 -0,556
 433 : begin twid_im = 32'b10010110011100111101101110010101; twid_re = 32'b10110111100101100001100110011100; end  //-0,825 -0,566
 434 : begin twid_im = 32'b10010111010110010110000110000000; twid_re = 32'b10110110010010111110101011001101; end  //-0,818 -0,576
 435 : begin twid_im = 32'b10011000010000101111000001000100; twid_re = 32'b10110101000001001001001101101001; end  //-0,810 -0,586
 436 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b10110011110000000010000000001101; end  //-0,803 -0,596
 437 : begin twid_im = 32'b10011010001000100000010000101110; twid_re = 32'b10110010011111101001110100111101; end  //-0,796 -0,606
 438 : begin twid_im = 32'b10011011000101110111011011011011; twid_re = 32'b10110001010000000001011101011100; end  //-0,788 -0,615
 439 : begin twid_im = 32'b10011100000100001100110101110001; twid_re = 32'b10110000000001001001101010110100; end  //-0,781 -0,625
 440 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b10101110110011000011001101101100; end  //-0,773 -0,634
 441 : begin twid_im = 32'b10011110000011101111111111000010; twid_re = 32'b10101101100101101110110110010010; end  //-0,765 -0,644
 442 : begin twid_im = 32'b10011111000100111100011111010001; twid_re = 32'b10101100011001001101010100010001; end  //-0,757 -0,653
 443 : begin twid_im = 32'b10100000000111000100110001110011; twid_re = 32'b10101011001101011111010110110110; end  //-0,749 -0,662
 444 : begin twid_im = 32'b10100001001010001000001101110111; twid_re = 32'b10101010000010100101101100101110; end  //-0,741 -0,672
 445 : begin twid_im = 32'b10100010001110000110001010000101; twid_re = 32'b10101000111000100001000100000111; end  //-0,733 -0,681
 446 : begin twid_im = 32'b10100011010010111101111100100001; twid_re = 32'b10100111101111010010001010101100; end  //-0,724 -0,690
 447 : begin twid_im = 32'b10100100011000101110111010101101; twid_re = 32'b10100110100110111001101101101001; end  //-0,716 -0,698
 448 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
 449 : begin twid_im = 32'b10100110100110111001101101101001; twid_re = 32'b10100100011000101110111010101101; end  //-0,698 -0,716
 450 : begin twid_im = 32'b10100111101111010010001010101100; twid_re = 32'b10100011010010111101111100100001; end  //-0,690 -0,724
 451 : begin twid_im = 32'b10101000111000100001000100000111; twid_re = 32'b10100010001110000110001010000101; end  //-0,681 -0,733
 452 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b10100001001010001000001101110111; end  //-0,672 -0,741
 453 : begin twid_im = 32'b10101011001101011111010110110110; twid_re = 32'b10100000000111000100110001110011; end  //-0,662 -0,749
 454 : begin twid_im = 32'b10101100011001001101010100010001; twid_re = 32'b10011111000100111100011111010001; end  //-0,653 -0,757
 455 : begin twid_im = 32'b10101101100101101110110110010010; twid_re = 32'b10011110000011101111111111000010; end  //-0,644 -0,765
 456 : begin twid_im = 32'b10101110110011000011001101101100; twid_re = 32'b10011101000011011111111001010100; end  //-0,634 -0,773
 457 : begin twid_im = 32'b10110000000001001001101010110100; twid_re = 32'b10011100000100001100110101110001; end  //-0,625 -0,781
 458 : begin twid_im = 32'b10110001010000000001011101011100; twid_re = 32'b10011011000101110111011011011011; end  //-0,615 -0,788
 459 : begin twid_im = 32'b10110010011111101001110100111101; twid_re = 32'b10011010001000100000010000101110; end  //-0,606 -0,796
 460 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b10011001001100000111111011100001; end  //-0,596 -0,803
 461 : begin twid_im = 32'b10110101000001001001001101101001; twid_re = 32'b10011000010000101111000001000100; end  //-0,586 -0,810
 462 : begin twid_im = 32'b10110110010010111110101011001101; twid_re = 32'b10010111010110010110000110000000; end  //-0,576 -0,818
 463 : begin twid_im = 32'b10110111100101100001100110011100; twid_re = 32'b10010110011100111101101110010101; end  //-0,566 -0,825
 464 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b10010101100100100110011101011101; end  //-0,556 -0,831
 465 : begin twid_im = 32'b10111010001100101100101001110001; twid_re = 32'b10010100101101010000110110001000; end  //-0,545 -0,838
 466 : begin twid_im = 32'b10111011100001010011001010110000; twid_re = 32'b10010011110110111101011010100001; end  //-0,535 -0,845
 467 : begin twid_im = 32'b10111100110110100011111011001011; twid_re = 32'b10010011000001101100101100000101; end  //-0,525 -0,851
 468 : begin twid_im = 32'b10111110001100011110000110011100; twid_re = 32'b10010010001101011111001011101100; end  //-0,514 -0,858
 469 : begin twid_im = 32'b10111111100011000000110111100011; twid_re = 32'b10010001011010010101011001100100; end  //-0,504 -0,864
 470 : begin twid_im = 32'b11000000111010001011011001001001; twid_re = 32'b10010000101000001111110101001111; end  //-0,493 -0,870
 471 : begin twid_im = 32'b11000010010001111100110101011011; twid_re = 32'b10001111110111001110111101100111; end  //-0,482 -0,876
 472 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b10001111000111010011010000111011; end  //-0,471 -0,882
 473 : begin twid_im = 32'b11000101000011010001000101001001; twid_re = 32'b10001110011000011101001100101111; end  //-0,461 -0,888
 474 : begin twid_im = 32'b11000110011100110010001011001110; twid_re = 32'b10001101101010101101001101111100; end  //-0,450 -0,893
 475 : begin twid_im = 32'b11000111110110110110110001010000; twid_re = 32'b10001100111110000011110000110001; end  //-0,439 -0,899
 476 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b10001100010010100001010000110000; end  //-0,428 -0,904
 477 : begin twid_im = 32'b11001010101100100110111110101010; twid_re = 32'b10001011101000000110001000110000; end  //-0,416 -0,909
 478 : begin twid_im = 32'b11001100001000010000110101111001; twid_re = 32'b10001010111110110010110010111100; end  //-0,405 -0,914
 479 : begin twid_im = 32'b11001101100100011010101100111001; twid_re = 32'b10001010010110100111101000110010; end  //-0,394 -0,919
 480 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b10001001101111100101000011000100; end  //-0,383 -0,924
 481 : begin twid_im = 32'b11010000011110001010110110011110; twid_re = 32'b10001001001001101011011001111000; end  //-0,371 -0,929
 482 : begin twid_im = 32'b11010001111011101111010110011110; twid_re = 32'b10001000100100111011000100100110; end  //-0,360 -0,933
 483 : begin twid_im = 32'b11010011011001110000010001000110; twid_re = 32'b10001000000001010100011001111000; end  //-0,348 -0,937
 484 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b10000111011110110111101111101101; end  //-0,337 -0,942
 485 : begin twid_im = 32'b11010110010111000011101101111011; twid_re = 32'b10000110111101100101011011010100; end  //-0,325 -0,946
 486 : begin twid_im = 32'b11010111110110010100011011011000; twid_re = 32'b10000110011101011101110001010000; end  //-0,314 -0,950
 487 : begin twid_im = 32'b11011001010101111101111001111011; twid_re = 32'b10000101111110100001000101010100; end  //-0,302 -0,953
 488 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b10000101100000101111101010100110; end  //-0,290 -0,957
 489 : begin twid_im = 32'b11011100010110010111011110000010; twid_re = 32'b10000101000100001001110011011101; end  //-0,279 -0,960
 490 : begin twid_im = 32'b11011101110111000101101100111011; twid_re = 32'b10000100101000101111110001100011; end  //-0,267 -0,964
 491 : begin twid_im = 32'b11011111011000001000111111100100; twid_re = 32'b10000100001110100001110101110001; end  //-0,255 -0,967
 492 : begin twid_im = 32'b11100000111001100000011010000101; twid_re = 32'b10000011110101100000010000010011; end  //-0,243 -0,970
 493 : begin twid_im = 32'b11100010011011001011000000011011; twid_re = 32'b10000011011101101011010000100011; end  //-0,231 -0,973
 494 : begin twid_im = 32'b11100011111101000111110110010110; twid_re = 32'b10000011000111000011000101001111; end  //-0,219 -0,976
 495 : begin twid_im = 32'b11100101011111010101111111011011; twid_re = 32'b10000010110001100111111100010101; end  //-0,207 -0,978
 496 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b10000010011101011010000011000001; end  //-0,195 -0,981
 497 : begin twid_im = 32'b11101000100100100010011000100010; twid_re = 32'b10000010001010011001100101110010; end  //-0,183 -0,983
 498 : begin twid_im = 32'b11101010000111011110101110111100; twid_re = 32'b10000001111000100110110000010111; end  //-0,171 -0,985
 499 : begin twid_im = 32'b11101011101010101000100101001111; twid_re = 32'b10000001101000000001101101101110; end  //-0,159 -0,987
 500 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b10000001011000101010101000000101; end  //-0,147 -0,989
 501 : begin twid_im = 32'b11101110110001100000111100110001; twid_re = 32'b10000001001010100001101000111011; end  //-0,135 -0,991
 502 : begin twid_im = 32'b11110000010101001101100011010101; twid_re = 32'b10000000111101100110111000111101; end  //-0,122 -0,992
 503 : begin twid_im = 32'b11110001111001000011110100011100; twid_re = 32'b10000000110001111010100000001011; end  //-0,110 -0,994
 504 : begin twid_im = 32'b11110011011101000010110010100010; twid_re = 32'b10000000100111011100100101110010; end  //-0,098 -0,995
 505 : begin twid_im = 32'b11110101000001001001011111111011; twid_re = 32'b10000000011110001101010000001110; end  //-0,086 -0,996
 506 : begin twid_im = 32'b11110110100101010110111110110111; twid_re = 32'b10000000010110001100100101001101; end  //-0,074 -0,997
 507 : begin twid_im = 32'b11111000001001101010010001100010; twid_re = 32'b10000000001111011010101001101011; end  //-0,061 -0,998
 508 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b10000000001001110111100001110011; end  //-0,049 -0,999
 509 : begin twid_im = 32'b11111011010010011110011010100011; twid_re = 32'b10000000000101100011010001000001; end  //-0,037 -0,999
 510 : begin twid_im = 32'b11111100110110111101010101000001; twid_re = 32'b10000000000010011101111001111111; end  //-0,025 -1,000
 511 : begin twid_im = 32'b11111110011011011110001011100000; twid_re = 32'b10000000000000100111011110100111; end  //-0,012 -1,000
 512 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 513 : begin twid_im = 32'b11111111001101101111000001111000; twid_re = 32'b01111111111111110110001000010101; end  //-0,006  1,000
 514 : begin twid_im = 32'b11111110011011011110001011100000; twid_re = 32'b01111111111111011000100001011001; end  //-0,012  1,000
 515 : begin twid_im = 32'b11111101101001001101100100101001; twid_re = 32'b01111111111110100111001011010000; end  //-0,018  1,000
 516 : begin twid_im = 32'b11111100110110111101010101000001; twid_re = 32'b01111111111101100010000110000001; end  //-0,025  1,000
 517 : begin twid_im = 32'b11111100000100101101100100011010; twid_re = 32'b01111111111100001001010001110111; end  //-0,031  1,000
 518 : begin twid_im = 32'b11111011010010011110011010100011; twid_re = 32'b01111111111010011100101110111111; end  //-0,037  0,999
 519 : begin twid_im = 32'b11111010100000001111111111001011; twid_re = 32'b01111111111000011100011101101010; end  //-0,043  0,999
 520 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b01111111110110001000011110001101; end  //-0,049  0,999
 521 : begin twid_im = 32'b11111000111011110101110010111011; twid_re = 32'b01111111110011100000110000111101; end  //-0,055  0,998
 522 : begin twid_im = 32'b11111000001001101010010001100010; twid_re = 32'b01111111110000100101010110010101; end  //-0,061  0,998
 523 : begin twid_im = 32'b11110111010111011111111101100110; twid_re = 32'b01111111101101010110001110110010; end  //-0,067  0,998
 524 : begin twid_im = 32'b11110110100101010110111110110111; twid_re = 32'b01111111101001110011011010110011; end  //-0,074  0,997
 525 : begin twid_im = 32'b11110101110011001111011101000100; twid_re = 32'b01111111100101111100111010111100; end  //-0,080  0,997
 526 : begin twid_im = 32'b11110101000001001001011111111011; twid_re = 32'b01111111100001110010101111110010; end  //-0,086  0,996
 527 : begin twid_im = 32'b11110100001111000101001111001011; twid_re = 32'b01111111011101010100111001111111; end  //-0,092  0,996
 528 : begin twid_im = 32'b11110011011101000010110010100010; twid_re = 32'b01111111011000100011011010001110; end  //-0,098  0,995
 529 : begin twid_im = 32'b11110010101011000010010001101110; twid_re = 32'b01111111010011011110010001010000; end  //-0,104  0,995
 530 : begin twid_im = 32'b11110001111001000011110100011100; twid_re = 32'b01111111001110000101011111110101; end  //-0,110  0,994
 531 : begin twid_im = 32'b11110001000111000111100010011010; twid_re = 32'b01111111001000011001000110110011; end  //-0,116  0,993
 532 : begin twid_im = 32'b11110000010101001101100011010101; twid_re = 32'b01111111000010011001000111000011; end  //-0,122  0,992
 533 : begin twid_im = 32'b11101111100011010101111110111000; twid_re = 32'b01111110111100000101100001011111; end  //-0,128  0,992
 534 : begin twid_im = 32'b11101110110001100000111100110001; twid_re = 32'b01111110110101011110010111000101; end  //-0,135  0,991
 535 : begin twid_im = 32'b11101101111111101110100100101011; twid_re = 32'b01111110101110100011101000111000; end  //-0,141  0,990
 536 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b01111110100111010101010111111011; end  //-0,147  0,989
 537 : begin twid_im = 32'b11101100011100010010010001001111; twid_re = 32'b01111110011111110011100101010110; end  //-0,153  0,988
 538 : begin twid_im = 32'b11101011101010101000100101001111; twid_re = 32'b01111110010111111110010010010010; end  //-0,159  0,987
 539 : begin twid_im = 32'b11101010111001000010000001111011; twid_re = 32'b01111110001111110101011111111110; end  //-0,165  0,986
 540 : begin twid_im = 32'b11101010000111011110101110111100; twid_re = 32'b01111110000111011001001111101001; end  //-0,171  0,985
 541 : begin twid_im = 32'b11101001010101111110110011111011; twid_re = 32'b01111101111110101001100010100111; end  //-0,177  0,984
 542 : begin twid_im = 32'b11101000100100100010011000100010; twid_re = 32'b01111101110101100110011010001110; end  //-0,183  0,983
 543 : begin twid_im = 32'b11100111110011001001100100011000; twid_re = 32'b01111101101100001111110111110111; end  //-0,189  0,982
 544 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b01111101100010100101111100111111; end  //-0,195  0,981
 545 : begin twid_im = 32'b11100110010000100011010000001101; twid_re = 32'b01111101011000101000101011000101; end  //-0,201  0,980
 546 : begin twid_im = 32'b11100101011111010101111111011011; twid_re = 32'b01111101001110011000000011101011; end  //-0,207  0,978
 547 : begin twid_im = 32'b11100100101110001100110100010001; twid_re = 32'b01111101000011110100001000010111; end  //-0,213  0,977
 548 : begin twid_im = 32'b11100011111101000111110110010110; twid_re = 32'b01111100111000111100111010110001; end  //-0,219  0,976
 549 : begin twid_im = 32'b11100011001100000111001101001101; twid_re = 32'b01111100101101110010011100100011; end  //-0,225  0,974
 550 : begin twid_im = 32'b11100010011011001011000000011011; twid_re = 32'b01111100100010010100101111011101; end  //-0,231  0,973
 551 : begin twid_im = 32'b11100001101010010011010111100010; twid_re = 32'b01111100010110100011110101001111; end  //-0,237  0,972
 552 : begin twid_im = 32'b11100000111001100000011010000101; twid_re = 32'b01111100001010011111101111101101; end  //-0,243  0,970
 553 : begin twid_im = 32'b11100000001000110010001111100101; twid_re = 32'b01111011111110001000100000101111; end  //-0,249  0,969
 554 : begin twid_im = 32'b11011111011000001000111111100100; twid_re = 32'b01111011110001011110001010001111; end  //-0,255  0,967
 555 : begin twid_im = 32'b11011110100111100100110001100001; twid_re = 32'b01111011100100100000101110001000; end  //-0,261  0,965
 556 : begin twid_im = 32'b11011101110111000101101100111011; twid_re = 32'b01111011010111010000001110011101; end  //-0,267  0,964
 557 : begin twid_im = 32'b11011101000110101011111001010001; twid_re = 32'b01111011001001101100101101001110; end  //-0,273  0,962
 558 : begin twid_im = 32'b11011100010110010111011110000010; twid_re = 32'b01111010111011110110001100100011; end  //-0,279  0,960
 559 : begin twid_im = 32'b11011011100110001000100010101001; twid_re = 32'b01111010101101101100101110100011; end  //-0,284  0,959
 560 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
 561 : begin twid_im = 32'b11011010000101111011101001001010; twid_re = 32'b01111010010000100001000011011000; end  //-0,296  0,955
 562 : begin twid_im = 32'b11011001010101111101111001111011; twid_re = 32'b01111010000001011110111010101100; end  //-0,302  0,953
 563 : begin twid_im = 32'b11011000100110000110001000001100; twid_re = 32'b01111001110010001001111101101101; end  //-0,308  0,951
 564 : begin twid_im = 32'b11010111110110010100011011011000; twid_re = 32'b01111001100010100010001110110000; end  //-0,314  0,950
 565 : begin twid_im = 32'b11010111000110101000111010110110; twid_re = 32'b01111001010010100111110000010001; end  //-0,320  0,948
 566 : begin twid_im = 32'b11010110010111000011101101111011; twid_re = 32'b01111001000010011010100100101100; end  //-0,325  0,946
 567 : begin twid_im = 32'b11010101100111100100111011111111; twid_re = 32'b01111000110001111010101110100001; end  //-0,331  0,944
 568 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b01111000100001001000010000010011; end  //-0,337  0,942
 569 : begin twid_im = 32'b11010100001000111011000110010001; twid_re = 32'b01111000010000000011001100101000; end  //-0,343  0,939
 570 : begin twid_im = 32'b11010011011001110000010001000110; twid_re = 32'b01110111111110101011100110001000; end  //-0,348  0,937
 571 : begin twid_im = 32'b11010010101010101100010100000101; twid_re = 32'b01110111101101000001011111011111; end  //-0,354  0,935
 572 : begin twid_im = 32'b11010001111011101111010110011110; twid_re = 32'b01110111011011000100111011011010; end  //-0,360  0,933
 573 : begin twid_im = 32'b11010001001100111001011111100010; twid_re = 32'b01110111001000110101111100101100; end  //-0,366  0,931
 574 : begin twid_im = 32'b11010000011110001010110110011110; twid_re = 32'b01110110110110010100100110001000; end  //-0,371  0,929
 575 : begin twid_im = 32'b11001111101111100011100010100000; twid_re = 32'b01110110100011100000111010100101; end  //-0,377  0,926
 576 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b01110110010000011010111100111100; end  //-0,383  0,924
 577 : begin twid_im = 32'b11001110010010101011010110100011; twid_re = 32'b01110101111101000010110000001010; end  //-0,388  0,922
 578 : begin twid_im = 32'b11001101100100011010101100111001; twid_re = 32'b01110101101001011000010111001110; end  //-0,394  0,919
 579 : begin twid_im = 32'b11001100110110010001110100111110; twid_re = 32'b01110101010101011011110101001011; end  //-0,400  0,917
 580 : begin twid_im = 32'b11001100001000010000110101111001; twid_re = 32'b01110101000001001101001101000100; end  //-0,405  0,914
 581 : begin twid_im = 32'b11001011011010010111110110110001; twid_re = 32'b01110100101100101100100010000011; end  //-0,411  0,912
 582 : begin twid_im = 32'b11001010101100100110111110101010; twid_re = 32'b01110100010111111001110111010000; end  //-0,416  0,909
 583 : begin twid_im = 32'b11001001111110111110010100100111; twid_re = 32'b01110100000010110101001111111010; end  //-0,422  0,907
 584 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b01110011101101011110101111010000; end  //-0,428  0,904
 585 : begin twid_im = 32'b11001000100100000110000110111010; twid_re = 32'b01110011010111110110011000100101; end  //-0,433  0,901
 586 : begin twid_im = 32'b11000111110110110110110001010000; twid_re = 32'b01110011000001111100001111001111; end  //-0,439  0,899
 587 : begin twid_im = 32'b11000111001001110000000101101101; twid_re = 32'b01110010101011110000010110100110; end  //-0,444  0,896
 588 : begin twid_im = 32'b11000110011100110010001011001110; twid_re = 32'b01110010010101010010110010000100; end  //-0,450  0,893
 589 : begin twid_im = 32'b11000101101111111101001000101111; twid_re = 32'b01110001111110100011100101001000; end  //-0,455  0,890
 590 : begin twid_im = 32'b11000101000011010001000101001001; twid_re = 32'b01110001100111100010110011010001; end  //-0,461  0,888
 591 : begin twid_im = 32'b11000100010110101110000111010111; twid_re = 32'b01110001010000010000100000000100; end  //-0,466  0,885
 592 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b01110000111000101100101111000101; end  //-0,471  0,882
 593 : begin twid_im = 32'b11000010111110000011111000101011; twid_re = 32'b01110000100000110111100011111110; end  //-0,477  0,879
 594 : begin twid_im = 32'b11000010010001111100110101011011; twid_re = 32'b01110000001000110001000010011001; end  //-0,482  0,876
 595 : begin twid_im = 32'b11000001100101111111010011010100; twid_re = 32'b01101111110000011001001110000100; end  //-0,488  0,873
 596 : begin twid_im = 32'b11000000111010001011011001001001; twid_re = 32'b01101111010111110000001010110001; end  //-0,493  0,870
 597 : begin twid_im = 32'b11000000001110100001001101101001; twid_re = 32'b01101110111110110101111100010001; end  //-0,498  0,867
 598 : begin twid_im = 32'b10111111100011000000110111100011; twid_re = 32'b01101110100101101010100110011100; end  //-0,504  0,864
 599 : begin twid_im = 32'b10111110110111101010011101100110; twid_re = 32'b01101110001100001110001101001001; end  //-0,509  0,861
 600 : begin twid_im = 32'b10111110001100011110000110011100; twid_re = 32'b01101101110010100000110100010100; end  //-0,514  0,858
 601 : begin twid_im = 32'b10111101100001011011111000110000; twid_re = 32'b01101101011000100010011111111001; end  //-0,519  0,855
 602 : begin twid_im = 32'b10111100110110100011111011001011; twid_re = 32'b01101100111110010011010011111011; end  //-0,525  0,851
 603 : begin twid_im = 32'b10111100001011110110010100010100; twid_re = 32'b01101100100011110011010100011011; end  //-0,530  0,848
 604 : begin twid_im = 32'b10111011100001010011001010110000; twid_re = 32'b01101100001001000010100101011111; end  //-0,535  0,845
 605 : begin twid_im = 32'b10111010110110111010100101000100; twid_re = 32'b01101011101110000001001011010000; end  //-0,540  0,842
 606 : begin twid_im = 32'b10111010001100101100101001110001; twid_re = 32'b01101011010010101111001001111000; end  //-0,545  0,838
 607 : begin twid_im = 32'b10111001100010101001011111011001; twid_re = 32'b01101010110111001100100101100100; end  //-0,550  0,835
 608 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
 609 : begin twid_im = 32'b10111000001111000011110111010010; twid_re = 32'b01101001111111010110000101001010; end  //-0,561  0,828
 610 : begin twid_im = 32'b10110111100101100001100110011100; twid_re = 32'b01101001100011000010010001101011; end  //-0,566  0,825
 611 : begin twid_im = 32'b10110110111100001010100000010010; twid_re = 32'b01101001000110011110001100011111; end  //-0,571  0,821
 612 : begin twid_im = 32'b10110110010010111110101011001101; twid_re = 32'b01101000101001101001111010000000; end  //-0,576  0,818
 613 : begin twid_im = 32'b10110101101001111110001101100011; twid_re = 32'b01101000001100100101011110101010; end  //-0,581  0,814
 614 : begin twid_im = 32'b10110101000001001001001101101001; twid_re = 32'b01100111101111010000111110111100; end  //-0,586  0,810
 615 : begin twid_im = 32'b10110100011000011111110001110001; twid_re = 32'b01100111010001101100011111010111; end  //-0,591  0,807
 616 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b01100110110011111000000100011111; end  //-0,596  0,803
 617 : begin twid_im = 32'b10110011000111101111111111001100; twid_re = 32'b01100110010101110011110010111011; end  //-0,601  0,800
 618 : begin twid_im = 32'b10110010011111101001110100111101; twid_re = 32'b01100101110111011111101111010010; end  //-0,606  0,796
 619 : begin twid_im = 32'b10110001110111101111100111101001; twid_re = 32'b01100101011000111011111110010001; end  //-0,610  0,792
 620 : begin twid_im = 32'b10110001010000000001011101011100; twid_re = 32'b01100100111010001000100100100101; end  //-0,615  0,788
 621 : begin twid_im = 32'b10110000101000011111011100011110; twid_re = 32'b01100100011011000101100110111111; end  //-0,620  0,785
 622 : begin twid_im = 32'b10110000000001001001101010110100; twid_re = 32'b01100011111011110011001010001111; end  //-0,625  0,781
 623 : begin twid_im = 32'b10101111011010000000001110100010; twid_re = 32'b01100011011100010001010011001100; end  //-0,630  0,777
 624 : begin twid_im = 32'b10101110110011000011001101101100; twid_re = 32'b01100010111100100000000110101100; end  //-0,634  0,773
 625 : begin twid_im = 32'b10101110001100010010101110010010; twid_re = 32'b01100010011100011111101001101000; end  //-0,639  0,769
 626 : begin twid_im = 32'b10101101100101101110110110010010; twid_re = 32'b01100001111100010000000000111110; end  //-0,644  0,765
 627 : begin twid_im = 32'b10101100111111010111101011101001; twid_re = 32'b01100001011011110001010001101011; end  //-0,649  0,761
 628 : begin twid_im = 32'b10101100011001001101010100010001; twid_re = 32'b01100000111011000011100000101111; end  //-0,653  0,757
 629 : begin twid_im = 32'b10101011110011001111110110000011; twid_re = 32'b01100000011010000110110011001110; end  //-0,658  0,753
 630 : begin twid_im = 32'b10101011001101011111010110110110; twid_re = 32'b01011111111000111011001110001101; end  //-0,662  0,749
 631 : begin twid_im = 32'b10101010100111111011111100011110; twid_re = 32'b01011111010111100000110110110010; end  //-0,667  0,745
 632 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b01011110110101110111110010001001; end  //-0,672  0,741
 633 : begin twid_im = 32'b10101001011101011100101101010111; twid_re = 32'b01011110010100000000000101011101; end  //-0,676  0,737
 634 : begin twid_im = 32'b10101000111000100001000100000111; twid_re = 32'b01011101110001111001110101111011; end  //-0,681  0,733
 635 : begin twid_im = 32'b10101000010011110010110110101011; twid_re = 32'b01011101001111100101001000110110; end  //-0,685  0,728
 636 : begin twid_im = 32'b10100111101111010010001010101100; twid_re = 32'b01011100101101000010000011011111; end  //-0,690  0,724
 637 : begin twid_im = 32'b10100111001010111111000101110100; twid_re = 32'b01011100001010010000101011001100; end  //-0,694  0,720
 638 : begin twid_im = 32'b10100110100110111001101101101001; twid_re = 32'b01011011100111010001000101010011; end  //-0,698  0,716
 639 : begin twid_im = 32'b10100110000011000010000111101110; twid_re = 32'b01011011000100000011010111001110; end  //-0,703  0,711
 640 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
 641 : begin twid_im = 32'b10100100111011111100101000110010; twid_re = 32'b01011001111100111101111000010010; end  //-0,711  0,703
 642 : begin twid_im = 32'b10100100011000101110111010101101; twid_re = 32'b01011001011001000110010010010111; end  //-0,716  0,698
 643 : begin twid_im = 32'b10100011110101101111010100110100; twid_re = 32'b01011000110101000000111010001100; end  //-0,720  0,694
 644 : begin twid_im = 32'b10100011010010111101111100100001; twid_re = 32'b01011000010000101101110101010100; end  //-0,724  0,690
 645 : begin twid_im = 32'b10100010110000011010110111001010; twid_re = 32'b01010111101100001101001001010101; end  //-0,728  0,685
 646 : begin twid_im = 32'b10100010001110000110001010000101; twid_re = 32'b01010111000111011110111011111001; end  //-0,733  0,681
 647 : begin twid_im = 32'b10100001101011111111111010100011; twid_re = 32'b01010110100010100011010010101001; end  //-0,737  0,676
 648 : begin twid_im = 32'b10100001001010001000001101110111; twid_re = 32'b01010101111101011010010011010010; end  //-0,741  0,672
 649 : begin twid_im = 32'b10100000101000011111001001001110; twid_re = 32'b01010101011000000100000011100010; end  //-0,745  0,667
 650 : begin twid_im = 32'b10100000000111000100110001110011; twid_re = 32'b01010100110010100000101001001010; end  //-0,749  0,662
 651 : begin twid_im = 32'b10011111100101111001001100110010; twid_re = 32'b01010100001100110000001001111101; end  //-0,753  0,658
 652 : begin twid_im = 32'b10011111000100111100011111010001; twid_re = 32'b01010011100110110010101011101111; end  //-0,757  0,653
 653 : begin twid_im = 32'b10011110100100001110101110010101; twid_re = 32'b01010011000000101000010100010111; end  //-0,761  0,649
 654 : begin twid_im = 32'b10011110000011101111111111000010; twid_re = 32'b01010010011010010001001001101110; end  //-0,765  0,644
 655 : begin twid_im = 32'b10011101100011100000010110011000; twid_re = 32'b01010001110011101101010001101110; end  //-0,769  0,639
 656 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
 657 : begin twid_im = 32'b10011100100011101110101100110100; twid_re = 32'b01010000100101111111110001011110; end  //-0,777  0,630
 658 : begin twid_im = 32'b10011100000100001100110101110001; twid_re = 32'b01001111111110110110010101001100; end  //-0,781  0,625
 659 : begin twid_im = 32'b10011011100100111010011001000001; twid_re = 32'b01001111010111100000100011100010; end  //-0,785  0,620
 660 : begin twid_im = 32'b10011011000101110111011011011011; twid_re = 32'b01001110101111111110100010100100; end  //-0,788  0,615
 661 : begin twid_im = 32'b10011010100111000100000001101111; twid_re = 32'b01001110001000010000011000010111; end  //-0,792  0,610
 662 : begin twid_im = 32'b10011010001000100000010000101110; twid_re = 32'b01001101100000010110001011000011; end  //-0,796  0,606
 663 : begin twid_im = 32'b10011001101010001100001101000101; twid_re = 32'b01001100111000010000000000110100; end  //-0,800  0,601
 664 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b01001100001111111101111111110011; end  //-0,803  0,596
 665 : begin twid_im = 32'b10011000101110010011100000101001; twid_re = 32'b01001011100111100000001110001111; end  //-0,807  0,591
 666 : begin twid_im = 32'b10011000010000101111000001000100; twid_re = 32'b01001010111110110110110010010111; end  //-0,810  0,586
 667 : begin twid_im = 32'b10010111110011011010100001010110; twid_re = 32'b01001010010110000001110010011101; end  //-0,814  0,581
 668 : begin twid_im = 32'b10010111010110010110000110000000; twid_re = 32'b01001001101101000001010100110011; end  //-0,818  0,576
 669 : begin twid_im = 32'b10010110111001100001110011100001; twid_re = 32'b01001001000011110101011111101110; end  //-0,821  0,571
 670 : begin twid_im = 32'b10010110011100111101101110010101; twid_re = 32'b01001000011010011110011001100100; end  //-0,825  0,566
 671 : begin twid_im = 32'b10010110000000101001111010110110; twid_re = 32'b01000111110000111100001000101110; end  //-0,828  0,561
 672 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b01000111000111001110110011100110; end  //-0,831  0,556
 673 : begin twid_im = 32'b10010101001000110011011010011100; twid_re = 32'b01000110011101010110100000100111; end  //-0,835  0,550
 674 : begin twid_im = 32'b10010100101101010000110110001000; twid_re = 32'b01000101110011010011010110001111; end  //-0,838  0,545
 675 : begin twid_im = 32'b10010100010001111110110100110000; twid_re = 32'b01000101001001000101011010111100; end  //-0,842  0,540
 676 : begin twid_im = 32'b10010011110110111101011010100001; twid_re = 32'b01000100011110101100110101010000; end  //-0,845  0,535
 677 : begin twid_im = 32'b10010011011100001100101011100101; twid_re = 32'b01000011110100001001101011101100; end  //-0,848  0,530
 678 : begin twid_im = 32'b10010011000001101100101100000101; twid_re = 32'b01000011001001011100000100110101; end  //-0,851  0,525
 679 : begin twid_im = 32'b10010010100111011101100000000111; twid_re = 32'b01000010011110100100000111010000; end  //-0,855  0,519
 680 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b01000001110011100001111001100100; end  //-0,858  0,514
 681 : begin twid_im = 32'b10010001110011110001110010110111; twid_re = 32'b01000001001000010101100010011010; end  //-0,861  0,509
 682 : begin twid_im = 32'b10010001011010010101011001100100; twid_re = 32'b01000000011100111111001000011101; end  //-0,864  0,504
 683 : begin twid_im = 32'b10010001000001001010000011101111; twid_re = 32'b00111111110001011110110010010111; end  //-0,867  0,498
 684 : begin twid_im = 32'b10010000101000001111110101001111; twid_re = 32'b00111111000101110100100110110111; end  //-0,870  0,493
 685 : begin twid_im = 32'b10010000001111100110110001111100; twid_re = 32'b00111110011010000000101100101100; end  //-0,873  0,488
 686 : begin twid_im = 32'b10001111110111001110111101100111; twid_re = 32'b00111101101110000011001010100101; end  //-0,876  0,482
 687 : begin twid_im = 32'b10001111011111001000011100000010; twid_re = 32'b00111101000001111100000111010101; end  //-0,879  0,477
 688 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b00111100010101101011101001110000; end  //-0,882  0,471
 689 : begin twid_im = 32'b10001110101111101111011111111100; twid_re = 32'b00111011101001010001111000101001; end  //-0,885  0,466
 690 : begin twid_im = 32'b10001110011000011101001100101111; twid_re = 32'b00111010111100101110111010110111; end  //-0,888  0,461
 691 : begin twid_im = 32'b10001110000001011100011010111000; twid_re = 32'b00111010010000000010110111010001; end  //-0,890  0,455
 692 : begin twid_im = 32'b10001101101010101101001101111100; twid_re = 32'b00111001100011001101110100110010; end  //-0,893  0,450
 693 : begin twid_im = 32'b10001101010100001111101001011010; twid_re = 32'b00111000110110001111111010010011; end  //-0,896  0,444
 694 : begin twid_im = 32'b10001100111110000011110000110001; twid_re = 32'b00111000001001001001001110110000; end  //-0,899  0,439
 695 : begin twid_im = 32'b10001100101000001001100111011011; twid_re = 32'b00110111011011111001111001000110; end  //-0,901  0,433
 696 : begin twid_im = 32'b10001100010010100001010000110000; twid_re = 32'b00110110101110100010000000010011; end  //-0,904  0,428
 697 : begin twid_im = 32'b10001011111101001010110000000110; twid_re = 32'b00110110000001000001101011011001; end  //-0,907  0,422
 698 : begin twid_im = 32'b10001011101000000110001000110000; twid_re = 32'b00110101010011011001000001010110; end  //-0,909  0,416
 699 : begin twid_im = 32'b10001011010011010011011101111101; twid_re = 32'b00110100100101101000001001001111; end  //-0,912  0,411
 700 : begin twid_im = 32'b10001010111110110010110010111100; twid_re = 32'b00110011110111101111001010000111; end  //-0,914  0,405
 701 : begin twid_im = 32'b10001010101010100100001010110101; twid_re = 32'b00110011001001101110001011000010; end  //-0,917  0,400
 702 : begin twid_im = 32'b10001010010110100111101000110010; twid_re = 32'b00110010011011100101010011000111; end  //-0,919  0,394
 703 : begin twid_im = 32'b10001010000010111101001111110110; twid_re = 32'b00110001101101010100101001011101; end  //-0,922  0,388
 704 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
 705 : begin twid_im = 32'b10001001011100011111000101011011; twid_re = 32'b00110000010000011100011101100000; end  //-0,926  0,377
 706 : begin twid_im = 32'b10001001001001101011011001111000; twid_re = 32'b00101111100001110101001001100010; end  //-0,929  0,371
 707 : begin twid_im = 32'b10001000110111001010000011010100; twid_re = 32'b00101110110011000110100000011110; end  //-0,931  0,366
 708 : begin twid_im = 32'b10001000100100111011000100100110; twid_re = 32'b00101110000100010000101001100010; end  //-0,933  0,360
 709 : begin twid_im = 32'b10001000010010111110100000100001; twid_re = 32'b00101101010101010011101011111011; end  //-0,935  0,354
 710 : begin twid_im = 32'b10001000000001010100011001111000; twid_re = 32'b00101100100110001111101110111010; end  //-0,937  0,348
 711 : begin twid_im = 32'b10000111101111111100110011011000; twid_re = 32'b00101011110111000100111001101111; end  //-0,939  0,343
 712 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b00101011000111110011010011101011; end  //-0,942  0,337
 713 : begin twid_im = 32'b10000111001110000101010001011111; twid_re = 32'b00101010011000011011000100000001; end  //-0,944  0,331
 714 : begin twid_im = 32'b10000110111101100101011011010100; twid_re = 32'b00101001101000111100010010000101; end  //-0,946  0,325
 715 : begin twid_im = 32'b10000110101101011000001111101111; twid_re = 32'b00101000111001010111000101001010; end  //-0,948  0,320
 716 : begin twid_im = 32'b10000110011101011101110001010000; twid_re = 32'b00101000001001101011100100101000; end  //-0,950  0,314
 717 : begin twid_im = 32'b10000110001101110110000010010011; twid_re = 32'b00100111011001111001110111110100; end  //-0,951  0,308
 718 : begin twid_im = 32'b10000101111110100001000101010100; twid_re = 32'b00100110101010000010000110000101; end  //-0,953  0,302
 719 : begin twid_im = 32'b10000101101111011110111100101000; twid_re = 32'b00100101111010000100010110110110; end  //-0,955  0,296
 720 : begin twid_im = 32'b10000101100000101111101010100110; twid_re = 32'b00100101001010000000110001011101; end  //-0,957  0,290
 721 : begin twid_im = 32'b10000101010010010011010001011101; twid_re = 32'b00100100011001110111011101010111; end  //-0,959  0,284
 722 : begin twid_im = 32'b10000101000100001001110011011101; twid_re = 32'b00100011101001101000100001111110; end  //-0,960  0,279
 723 : begin twid_im = 32'b10000100110110010011010010110010; twid_re = 32'b00100010111001010100000110101111; end  //-0,962  0,273
 724 : begin twid_im = 32'b10000100101000101111110001100011; twid_re = 32'b00100010001000111010010011000101; end  //-0,964  0,267
 725 : begin twid_im = 32'b10000100011011011111010001111000; twid_re = 32'b00100001011000011011001110011111; end  //-0,965  0,261
 726 : begin twid_im = 32'b10000100001110100001110101110001; twid_re = 32'b00100000100111110111000000011100; end  //-0,967  0,255
 727 : begin twid_im = 32'b10000100000001110111011111010001; twid_re = 32'b00011111110111001101110000011011; end  //-0,969  0,249
 728 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b00011111000110011111100101111011; end  //-0,970  0,243
 729 : begin twid_im = 32'b10000011101001011100001010110001; twid_re = 32'b00011110010101101100101000011110; end  //-0,972  0,237
 730 : begin twid_im = 32'b10000011011101101011010000100011; twid_re = 32'b00011101100100110100111111100101; end  //-0,973  0,231
 731 : begin twid_im = 32'b10000011010010001101100011011101; twid_re = 32'b00011100110011111000110010110011; end  //-0,974  0,225
 732 : begin twid_im = 32'b10000011000111000011000101001111; twid_re = 32'b00011100000010111000001001101010; end  //-0,976  0,219
 733 : begin twid_im = 32'b10000010111100001011110111101001; twid_re = 32'b00011011010001110011001011101111; end  //-0,977  0,213
 734 : begin twid_im = 32'b10000010110001100111111100010101; twid_re = 32'b00011010100000101010000000100101; end  //-0,978  0,207
 735 : begin twid_im = 32'b10000010100111010111010100111011; twid_re = 32'b00011001101111011100101111110011; end  //-0,980  0,201
 736 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b00011000111110001011100000111100; end  //-0,981  0,195
 737 : begin twid_im = 32'b10000010010011110000001000001001; twid_re = 32'b00011000001100110110011011101000; end  //-0,982  0,189
 738 : begin twid_im = 32'b10000010001010011001100101110010; twid_re = 32'b00010111011011011101100111011110; end  //-0,983  0,183
 739 : begin twid_im = 32'b10000010000001010110011101011001; twid_re = 32'b00010110101010000001001100000101; end  //-0,984  0,177
 740 : begin twid_im = 32'b10000001111000100110110000010111; twid_re = 32'b00010101111000100001010001000100; end  //-0,985  0,171
 741 : begin twid_im = 32'b10000001110000001010100000000010; twid_re = 32'b00010101000110111101111110000101; end  //-0,986  0,165
 742 : begin twid_im = 32'b10000001101000000001101101101110; twid_re = 32'b00010100010101010111011010110001; end  //-0,987  0,159
 743 : begin twid_im = 32'b10000001100000001100011010101010; twid_re = 32'b00010011100011101101101110110001; end  //-0,988  0,153
 744 : begin twid_im = 32'b10000001011000101010101000000101; twid_re = 32'b00010010110010000001000001101110; end  //-0,989  0,147
 745 : begin twid_im = 32'b10000001010001011100010111001000; twid_re = 32'b00010010000000010001011011010101; end  //-0,990  0,141
 746 : begin twid_im = 32'b10000001001010100001101000111011; twid_re = 32'b00010001001110011111000011001111; end  //-0,991  0,135
 747 : begin twid_im = 32'b10000001000011111010011110100001; twid_re = 32'b00010000011100101010000001001000; end  //-0,992  0,128
 748 : begin twid_im = 32'b10000000111101100110111000111101; twid_re = 32'b00001111101010110010011100101011; end  //-0,992  0,122
 749 : begin twid_im = 32'b10000000110111100110111001001101; twid_re = 32'b00001110111000111000011101100110; end  //-0,993  0,116
 750 : begin twid_im = 32'b10000000110001111010100000001011; twid_re = 32'b00001110000110111100001011100100; end  //-0,994  0,110
 751 : begin twid_im = 32'b10000000101100100001101110110000; twid_re = 32'b00001101010100111101101110010010; end  //-0,995  0,104
 752 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
 753 : begin twid_im = 32'b10000000100010101011000110000001; twid_re = 32'b00001011110000111010110000110101; end  //-0,996  0,092
 754 : begin twid_im = 32'b10000000011110001101010000001110; twid_re = 32'b00001010111110110110100000000101; end  //-0,996  0,086
 755 : begin twid_im = 32'b10000000011010000011000101000100; twid_re = 32'b00001010001100110000100010111100; end  //-0,997  0,080
 756 : begin twid_im = 32'b10000000010110001100100101001101; twid_re = 32'b00001001011010101001000001001001; end  //-0,997  0,074
 757 : begin twid_im = 32'b10000000010010101001110001001110; twid_re = 32'b00001000101000100000000010011010; end  //-0,998  0,067
 758 : begin twid_im = 32'b10000000001111011010101001101011; twid_re = 32'b00000111110110010101101110011110; end  //-0,998  0,061
 759 : begin twid_im = 32'b10000000001100011111001111000011; twid_re = 32'b00000111000100001010001101000101; end  //-0,998  0,055
 760 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b00000110010001111101100101111100; end  //-0,999  0,049
 761 : begin twid_im = 32'b10000000000111100011100010010110; twid_re = 32'b00000101011111110000000000110101; end  //-0,999  0,043
 762 : begin twid_im = 32'b10000000000101100011010001000001; twid_re = 32'b00000100101101100001100101011101; end  //-0,999  0,037
 763 : begin twid_im = 32'b10000000000011110110101110001001; twid_re = 32'b00000011111011010010011011100110; end  //-1,000  0,031
 764 : begin twid_im = 32'b10000000000010011101111001111111; twid_re = 32'b00000011001001000010101010111111; end  //-1,000  0,025
 765 : begin twid_im = 32'b10000000000001011000110100110000; twid_re = 32'b00000010010110110010011011010111; end  //-1,000  0,018
 766 : begin twid_im = 32'b10000000000000100111011110100111; twid_re = 32'b00000001100100100001110100100000; end  //-1,000  0,012
 767 : begin twid_im = 32'b10000000000000001001110111101011; twid_re = 32'b00000000110010010000111110001000; end  //-1,000  0,006
 768 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 769 : begin twid_im = 32'b11111101101001001101100100101001; twid_re = 32'b01111111111110100111001011010000; end  //-0,018  1,000
 770 : begin twid_im = 32'b11111011010010011110011010100011; twid_re = 32'b01111111111010011100101110111111; end  //-0,037  0,999
 771 : begin twid_im = 32'b11111000111011110101110010111011; twid_re = 32'b01111111110011100000110000111101; end  //-0,055  0,998
 772 : begin twid_im = 32'b11110110100101010110111110110111; twid_re = 32'b01111111101001110011011010110011; end  //-0,074  0,997
 773 : begin twid_im = 32'b11110100001111000101001111001011; twid_re = 32'b01111111011101010100111001111111; end  //-0,092  0,996
 774 : begin twid_im = 32'b11110001111001000011110100011100; twid_re = 32'b01111111001110000101011111110101; end  //-0,110  0,994
 775 : begin twid_im = 32'b11101111100011010101111110111000; twid_re = 32'b01111110111100000101100001011111; end  //-0,128  0,992
 776 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b01111110100111010101010111111011; end  //-0,147  0,989
 777 : begin twid_im = 32'b11101010111001000010000001111011; twid_re = 32'b01111110001111110101011111111110; end  //-0,165  0,986
 778 : begin twid_im = 32'b11101000100100100010011000100010; twid_re = 32'b01111101110101100110011010001110; end  //-0,183  0,983
 779 : begin twid_im = 32'b11100110010000100011010000001101; twid_re = 32'b01111101011000101000101011000101; end  //-0,201  0,980
 780 : begin twid_im = 32'b11100011111101000111110110010110; twid_re = 32'b01111100111000111100111010110001; end  //-0,219  0,976
 781 : begin twid_im = 32'b11100001101010010011010111100010; twid_re = 32'b01111100010110100011110101001111; end  //-0,237  0,972
 782 : begin twid_im = 32'b11011111011000001000111111100100; twid_re = 32'b01111011110001011110001010001111; end  //-0,255  0,967
 783 : begin twid_im = 32'b11011101000110101011111001010001; twid_re = 32'b01111011001001101100101101001110; end  //-0,273  0,962
 784 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
 785 : begin twid_im = 32'b11011000100110000110001000001100; twid_re = 32'b01111001110010001001111101101101; end  //-0,308  0,951
 786 : begin twid_im = 32'b11010110010111000011101101111011; twid_re = 32'b01111001000010011010100100101100; end  //-0,325  0,946
 787 : begin twid_im = 32'b11010100001000111011000110010001; twid_re = 32'b01111000010000000011001100101000; end  //-0,343  0,939
 788 : begin twid_im = 32'b11010001111011101111010110011110; twid_re = 32'b01110111011011000100111011011010; end  //-0,360  0,933
 789 : begin twid_im = 32'b11001111101111100011100010100000; twid_re = 32'b01110110100011100000111010100101; end  //-0,377  0,926
 790 : begin twid_im = 32'b11001101100100011010101100111001; twid_re = 32'b01110101101001011000010111001110; end  //-0,394  0,919
 791 : begin twid_im = 32'b11001011011010010111110110110001; twid_re = 32'b01110100101100101100100010000011; end  //-0,411  0,912
 792 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b01110011101101011110101111010000; end  //-0,428  0,904
 793 : begin twid_im = 32'b11000111001001110000000101101101; twid_re = 32'b01110010101011110000010110100110; end  //-0,444  0,896
 794 : begin twid_im = 32'b11000101000011010001000101001001; twid_re = 32'b01110001100111100010110011010001; end  //-0,461  0,888
 795 : begin twid_im = 32'b11000010111110000011111000101011; twid_re = 32'b01110000100000110111100011111110; end  //-0,477  0,879
 796 : begin twid_im = 32'b11000000111010001011011001001001; twid_re = 32'b01101111010111110000001010110001; end  //-0,493  0,870
 797 : begin twid_im = 32'b10111110110111101010011101100110; twid_re = 32'b01101110001100001110001101001001; end  //-0,509  0,861
 798 : begin twid_im = 32'b10111100110110100011111011001011; twid_re = 32'b01101100111110010011010011111011; end  //-0,525  0,851
 799 : begin twid_im = 32'b10111010110110111010100101000100; twid_re = 32'b01101011101110000001001011010000; end  //-0,540  0,842
 800 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
 801 : begin twid_im = 32'b10110110111100001010100000010010; twid_re = 32'b01101001000110011110001100011111; end  //-0,571  0,821
 802 : begin twid_im = 32'b10110101000001001001001101101001; twid_re = 32'b01100111101111010000111110111100; end  //-0,586  0,810
 803 : begin twid_im = 32'b10110011000111101111111111001100; twid_re = 32'b01100110010101110011110010111011; end  //-0,601  0,800
 804 : begin twid_im = 32'b10110001010000000001011101011100; twid_re = 32'b01100100111010001000100100100101; end  //-0,615  0,788
 805 : begin twid_im = 32'b10101111011010000000001110100010; twid_re = 32'b01100011011100010001010011001100; end  //-0,630  0,777
 806 : begin twid_im = 32'b10101101100101101110110110010010; twid_re = 32'b01100001111100010000000000111110; end  //-0,644  0,765
 807 : begin twid_im = 32'b10101011110011001111110110000011; twid_re = 32'b01100000011010000110110011001110; end  //-0,658  0,753
 808 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b01011110110101110111110010001001; end  //-0,672  0,741
 809 : begin twid_im = 32'b10101000010011110010110110101011; twid_re = 32'b01011101001111100101001000110110; end  //-0,685  0,728
 810 : begin twid_im = 32'b10100110100110111001101101101001; twid_re = 32'b01011011100111010001000101010011; end  //-0,698  0,716
 811 : begin twid_im = 32'b10100100111011111100101000110010; twid_re = 32'b01011001111100111101111000010010; end  //-0,711  0,703
 812 : begin twid_im = 32'b10100011010010111101111100100001; twid_re = 32'b01011000010000101101110101010100; end  //-0,724  0,690
 813 : begin twid_im = 32'b10100001101011111111111010100011; twid_re = 32'b01010110100010100011010010101001; end  //-0,737  0,676
 814 : begin twid_im = 32'b10100000000111000100110001110011; twid_re = 32'b01010100110010100000101001001010; end  //-0,749  0,662
 815 : begin twid_im = 32'b10011110100100001110101110010101; twid_re = 32'b01010011000000101000010100010111; end  //-0,761  0,649
 816 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
 817 : begin twid_im = 32'b10011011100100111010011001000001; twid_re = 32'b01001111010111100000100011100010; end  //-0,785  0,620
 818 : begin twid_im = 32'b10011010001000100000010000101110; twid_re = 32'b01001101100000010110001011000011; end  //-0,796  0,606
 819 : begin twid_im = 32'b10011000101110010011100000101001; twid_re = 32'b01001011100111100000001110001111; end  //-0,807  0,591
 820 : begin twid_im = 32'b10010111010110010110000110000000; twid_re = 32'b01001001101101000001010100110011; end  //-0,818  0,576
 821 : begin twid_im = 32'b10010110000000101001111010110110; twid_re = 32'b01000111110000111100001000101110; end  //-0,828  0,561
 822 : begin twid_im = 32'b10010100101101010000110110001000; twid_re = 32'b01000101110011010011010110001111; end  //-0,838  0,545
 823 : begin twid_im = 32'b10010011011100001100101011100101; twid_re = 32'b01000011110100001001101011101100; end  //-0,848  0,530
 824 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b01000001110011100001111001100100; end  //-0,858  0,514
 825 : begin twid_im = 32'b10010001000001001010000011101111; twid_re = 32'b00111111110001011110110010010111; end  //-0,867  0,498
 826 : begin twid_im = 32'b10001111110111001110111101100111; twid_re = 32'b00111101101110000011001010100101; end  //-0,876  0,482
 827 : begin twid_im = 32'b10001110101111101111011111111100; twid_re = 32'b00111011101001010001111000101001; end  //-0,885  0,466
 828 : begin twid_im = 32'b10001101101010101101001101111100; twid_re = 32'b00111001100011001101110100110010; end  //-0,893  0,450
 829 : begin twid_im = 32'b10001100101000001001100111011011; twid_re = 32'b00110111011011111001111001000110; end  //-0,901  0,433
 830 : begin twid_im = 32'b10001011101000000110001000110000; twid_re = 32'b00110101010011011001000001010110; end  //-0,909  0,416
 831 : begin twid_im = 32'b10001010101010100100001010110101; twid_re = 32'b00110011001001101110001011000010; end  //-0,917  0,400
 832 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
 833 : begin twid_im = 32'b10001000110111001010000011010100; twid_re = 32'b00101110110011000110100000011110; end  //-0,931  0,366
 834 : begin twid_im = 32'b10001000000001010100011001111000; twid_re = 32'b00101100100110001111101110111010; end  //-0,937  0,348
 835 : begin twid_im = 32'b10000111001110000101010001011111; twid_re = 32'b00101010011000011011000100000001; end  //-0,944  0,331
 836 : begin twid_im = 32'b10000110011101011101110001010000; twid_re = 32'b00101000001001101011100100101000; end  //-0,950  0,314
 837 : begin twid_im = 32'b10000101101111011110111100101000; twid_re = 32'b00100101111010000100010110110110; end  //-0,955  0,296
 838 : begin twid_im = 32'b10000101000100001001110011011101; twid_re = 32'b00100011101001101000100001111110; end  //-0,960  0,279
 839 : begin twid_im = 32'b10000100011011011111010001111000; twid_re = 32'b00100001011000011011001110011111; end  //-0,965  0,261
 840 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b00011111000110011111100101111011; end  //-0,970  0,243
 841 : begin twid_im = 32'b10000011010010001101100011011101; twid_re = 32'b00011100110011111000110010110011; end  //-0,974  0,225
 842 : begin twid_im = 32'b10000010110001100111111100010101; twid_re = 32'b00011010100000101010000000100101; end  //-0,978  0,207
 843 : begin twid_im = 32'b10000010010011110000001000001001; twid_re = 32'b00011000001100110110011011101000; end  //-0,982  0,189
 844 : begin twid_im = 32'b10000001111000100110110000010111; twid_re = 32'b00010101111000100001010001000100; end  //-0,985  0,171
 845 : begin twid_im = 32'b10000001100000001100011010101010; twid_re = 32'b00010011100011101101101110110001; end  //-0,988  0,153
 846 : begin twid_im = 32'b10000001001010100001101000111011; twid_re = 32'b00010001001110011111000011001111; end  //-0,991  0,135
 847 : begin twid_im = 32'b10000000110111100110111001001101; twid_re = 32'b00001110111000111000011101100110; end  //-0,993  0,116
 848 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
 849 : begin twid_im = 32'b10000000011010000011000101000100; twid_re = 32'b00001010001100110000100010111100; end  //-0,997  0,080
 850 : begin twid_im = 32'b10000000001111011010101001101011; twid_re = 32'b00000111110110010101101110011110; end  //-0,998  0,061
 851 : begin twid_im = 32'b10000000000111100011100010010110; twid_re = 32'b00000101011111110000000000110101; end  //-0,999  0,043
 852 : begin twid_im = 32'b10000000000010011101111001111111; twid_re = 32'b00000011001001000010101010111111; end  //-1,000  0,025
 853 : begin twid_im = 32'b10000000000000001001110111101011; twid_re = 32'b00000000110010010000111110001000; end  //-1,000  0,006
 854 : begin twid_im = 32'b10000000000000100111011110100111; twid_re = 32'b11111110011011011110001011100000; end  //-1,000 -0,012
 855 : begin twid_im = 32'b10000000000011110110101110001001; twid_re = 32'b11111100000100101101100100011010; end  //-1,000 -0,031
 856 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b11111001101110000010011010000100; end  //-0,999 -0,049
 857 : begin twid_im = 32'b10000000010010101001110001001110; twid_re = 32'b11110111010111011111111101100110; end  //-0,998 -0,067
 858 : begin twid_im = 32'b10000000011110001101010000001110; twid_re = 32'b11110101000001001001011111111011; end  //-0,996 -0,086
 859 : begin twid_im = 32'b10000000101100100001101110110000; twid_re = 32'b11110010101011000010010001101110; end  //-0,995 -0,104
 860 : begin twid_im = 32'b10000000111101100110111000111101; twid_re = 32'b11110000010101001101100011010101; end  //-0,992 -0,122
 861 : begin twid_im = 32'b10000001010001011100010111001000; twid_re = 32'b11101101111111101110100100101011; end  //-0,990 -0,141
 862 : begin twid_im = 32'b10000001101000000001101101101110; twid_re = 32'b11101011101010101000100101001111; end  //-0,987 -0,159
 863 : begin twid_im = 32'b10000010000001010110011101011001; twid_re = 32'b11101001010101111110110011111011; end  //-0,984 -0,177
 864 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b11100111000001110100011111000100; end  //-0,981 -0,195
 865 : begin twid_im = 32'b10000010111100001011110111101001; twid_re = 32'b11100100101110001100110100010001; end  //-0,977 -0,213
 866 : begin twid_im = 32'b10000011011101101011010000100011; twid_re = 32'b11100010011011001011000000011011; end  //-0,973 -0,231
 867 : begin twid_im = 32'b10000100000001110111011111010001; twid_re = 32'b11100000001000110010001111100101; end  //-0,969 -0,249
 868 : begin twid_im = 32'b10000100101000101111110001100011; twid_re = 32'b11011101110111000101101100111011; end  //-0,964 -0,267
 869 : begin twid_im = 32'b10000101010010010011010001011101; twid_re = 32'b11011011100110001000100010101001; end  //-0,959 -0,284
 870 : begin twid_im = 32'b10000101111110100001000101010100; twid_re = 32'b11011001010101111101111001111011; end  //-0,953 -0,302
 871 : begin twid_im = 32'b10000110101101011000001111101111; twid_re = 32'b11010111000110101000111010110110; end  //-0,948 -0,320
 872 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b11010100111000001100101100010101; end  //-0,942 -0,337
 873 : begin twid_im = 32'b10001000010010111110100000100001; twid_re = 32'b11010010101010101100010100000101; end  //-0,935 -0,354
 874 : begin twid_im = 32'b10001001001001101011011001111000; twid_re = 32'b11010000011110001010110110011110; end  //-0,929 -0,371
 875 : begin twid_im = 32'b10001010000010111101001111110110; twid_re = 32'b11001110010010101011010110100011; end  //-0,922 -0,388
 876 : begin twid_im = 32'b10001010111110110010110010111100; twid_re = 32'b11001100001000010000110101111001; end  //-0,914 -0,405
 877 : begin twid_im = 32'b10001011111101001010110000000110; twid_re = 32'b11001001111110111110010100100111; end  //-0,907 -0,422
 878 : begin twid_im = 32'b10001100111110000011110000110001; twid_re = 32'b11000111110110110110110001010000; end  //-0,899 -0,439
 879 : begin twid_im = 32'b10001110000001011100011010111000; twid_re = 32'b11000101101111111101001000101111; end  //-0,890 -0,455
 880 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b11000011101010010100010110010000; end  //-0,882 -0,471
 881 : begin twid_im = 32'b10010000001111100110110001111100; twid_re = 32'b11000001100101111111010011010100; end  //-0,873 -0,488
 882 : begin twid_im = 32'b10010001011010010101011001100100; twid_re = 32'b10111111100011000000110111100011; end  //-0,864 -0,504
 883 : begin twid_im = 32'b10010010100111011101100000000111; twid_re = 32'b10111101100001011011111000110000; end  //-0,855 -0,519
 884 : begin twid_im = 32'b10010011110110111101011010100001; twid_re = 32'b10111011100001010011001010110000; end  //-0,845 -0,535
 885 : begin twid_im = 32'b10010101001000110011011010011100; twid_re = 32'b10111001100010101001011111011001; end  //-0,835 -0,550
 886 : begin twid_im = 32'b10010110011100111101101110010101; twid_re = 32'b10110111100101100001100110011100; end  //-0,825 -0,566
 887 : begin twid_im = 32'b10010111110011011010100001010110; twid_re = 32'b10110101101001111110001101100011; end  //-0,814 -0,581
 888 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b10110011110000000010000000001101; end  //-0,803 -0,596
 889 : begin twid_im = 32'b10011010100111000100000001101111; twid_re = 32'b10110001110111101111100111101001; end  //-0,792 -0,610
 890 : begin twid_im = 32'b10011100000100001100110101110001; twid_re = 32'b10110000000001001001101010110100; end  //-0,781 -0,625
 891 : begin twid_im = 32'b10011101100011100000010110011000; twid_re = 32'b10101110001100010010101110010010; end  //-0,769 -0,639
 892 : begin twid_im = 32'b10011111000100111100011111010001; twid_re = 32'b10101100011001001101010100010001; end  //-0,757 -0,653
 893 : begin twid_im = 32'b10100000101000011111001001001110; twid_re = 32'b10101010100111111011111100011110; end  //-0,745 -0,667
 894 : begin twid_im = 32'b10100010001110000110001010000101; twid_re = 32'b10101000111000100001000100000111; end  //-0,733 -0,681
 895 : begin twid_im = 32'b10100011110101101111010100110100; twid_re = 32'b10100111001010111111000101110100; end  //-0,720 -0,694
 896 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
 897 : begin twid_im = 32'b10100111001010111111000101110100; twid_re = 32'b10100011110101101111010100110100; end  //-0,694 -0,720
 898 : begin twid_im = 32'b10101000111000100001000100000111; twid_re = 32'b10100010001110000110001010000101; end  //-0,681 -0,733
 899 : begin twid_im = 32'b10101010100111111011111100011110; twid_re = 32'b10100000101000011111001001001110; end  //-0,667 -0,745
 900 : begin twid_im = 32'b10101100011001001101010100010001; twid_re = 32'b10011111000100111100011111010001; end  //-0,653 -0,757
 901 : begin twid_im = 32'b10101110001100010010101110010010; twid_re = 32'b10011101100011100000010110011000; end  //-0,639 -0,769
 902 : begin twid_im = 32'b10110000000001001001101010110100; twid_re = 32'b10011100000100001100110101110001; end  //-0,625 -0,781
 903 : begin twid_im = 32'b10110001110111101111100111101001; twid_re = 32'b10011010100111000100000001101111; end  //-0,610 -0,792
 904 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b10011001001100000111111011100001; end  //-0,596 -0,803
 905 : begin twid_im = 32'b10110101101001111110001101100011; twid_re = 32'b10010111110011011010100001010110; end  //-0,581 -0,814
 906 : begin twid_im = 32'b10110111100101100001100110011100; twid_re = 32'b10010110011100111101101110010101; end  //-0,566 -0,825
 907 : begin twid_im = 32'b10111001100010101001011111011001; twid_re = 32'b10010101001000110011011010011100; end  //-0,550 -0,835
 908 : begin twid_im = 32'b10111011100001010011001010110000; twid_re = 32'b10010011110110111101011010100001; end  //-0,535 -0,845
 909 : begin twid_im = 32'b10111101100001011011111000110000; twid_re = 32'b10010010100111011101100000000111; end  //-0,519 -0,855
 910 : begin twid_im = 32'b10111111100011000000110111100011; twid_re = 32'b10010001011010010101011001100100; end  //-0,504 -0,864
 911 : begin twid_im = 32'b11000001100101111111010011010100; twid_re = 32'b10010000001111100110110001111100; end  //-0,488 -0,873
 912 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b10001111000111010011010000111011; end  //-0,471 -0,882
 913 : begin twid_im = 32'b11000101101111111101001000101111; twid_re = 32'b10001110000001011100011010111000; end  //-0,455 -0,890
 914 : begin twid_im = 32'b11000111110110110110110001010000; twid_re = 32'b10001100111110000011110000110001; end  //-0,439 -0,899
 915 : begin twid_im = 32'b11001001111110111110010100100111; twid_re = 32'b10001011111101001010110000000110; end  //-0,422 -0,907
 916 : begin twid_im = 32'b11001100001000010000110101111001; twid_re = 32'b10001010111110110010110010111100; end  //-0,405 -0,914
 917 : begin twid_im = 32'b11001110010010101011010110100011; twid_re = 32'b10001010000010111101001111110110; end  //-0,388 -0,922
 918 : begin twid_im = 32'b11010000011110001010110110011110; twid_re = 32'b10001001001001101011011001111000; end  //-0,371 -0,929
 919 : begin twid_im = 32'b11010010101010101100010100000101; twid_re = 32'b10001000010010111110100000100001; end  //-0,354 -0,935
 920 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b10000111011110110111101111101101; end  //-0,337 -0,942
 921 : begin twid_im = 32'b11010111000110101000111010110110; twid_re = 32'b10000110101101011000001111101111; end  //-0,320 -0,948
 922 : begin twid_im = 32'b11011001010101111101111001111011; twid_re = 32'b10000101111110100001000101010100; end  //-0,302 -0,953
 923 : begin twid_im = 32'b11011011100110001000100010101001; twid_re = 32'b10000101010010010011010001011101; end  //-0,284 -0,959
 924 : begin twid_im = 32'b11011101110111000101101100111011; twid_re = 32'b10000100101000101111110001100011; end  //-0,267 -0,964
 925 : begin twid_im = 32'b11100000001000110010001111100101; twid_re = 32'b10000100000001110111011111010001; end  //-0,249 -0,969
 926 : begin twid_im = 32'b11100010011011001011000000011011; twid_re = 32'b10000011011101101011010000100011; end  //-0,231 -0,973
 927 : begin twid_im = 32'b11100100101110001100110100010001; twid_re = 32'b10000010111100001011110111101001; end  //-0,213 -0,977
 928 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b10000010011101011010000011000001; end  //-0,195 -0,981
 929 : begin twid_im = 32'b11101001010101111110110011111011; twid_re = 32'b10000010000001010110011101011001; end  //-0,177 -0,984
 930 : begin twid_im = 32'b11101011101010101000100101001111; twid_re = 32'b10000001101000000001101101101110; end  //-0,159 -0,987
 931 : begin twid_im = 32'b11101101111111101110100100101011; twid_re = 32'b10000001010001011100010111001000; end  //-0,141 -0,990
 932 : begin twid_im = 32'b11110000010101001101100011010101; twid_re = 32'b10000000111101100110111000111101; end  //-0,122 -0,992
 933 : begin twid_im = 32'b11110010101011000010010001101110; twid_re = 32'b10000000101100100001101110110000; end  //-0,104 -0,995
 934 : begin twid_im = 32'b11110101000001001001011111111011; twid_re = 32'b10000000011110001101010000001110; end  //-0,086 -0,996
 935 : begin twid_im = 32'b11110111010111011111111101100110; twid_re = 32'b10000000010010101001110001001110; end  //-0,067 -0,998
 936 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b10000000001001110111100001110011; end  //-0,049 -0,999
 937 : begin twid_im = 32'b11111100000100101101100100011010; twid_re = 32'b10000000000011110110101110001001; end  //-0,031 -1,000
 938 : begin twid_im = 32'b11111110011011011110001011100000; twid_re = 32'b10000000000000100111011110100111; end  //-0,012 -1,000
 939 : begin twid_im = 32'b00000000110010010000111110001000; twid_re = 32'b10000000000000001001110111101011; end  // 0,006 -1,000
 940 : begin twid_im = 32'b00000011001001000010101010111111; twid_re = 32'b10000000000010011101111001111111; end  // 0,025 -1,000
 941 : begin twid_im = 32'b00000101011111110000000000110101; twid_re = 32'b10000000000111100011100010010110; end  // 0,043 -0,999
 942 : begin twid_im = 32'b00000111110110010101101110011110; twid_re = 32'b10000000001111011010101001101011; end  // 0,061 -0,998
 943 : begin twid_im = 32'b00001010001100110000100010111100; twid_re = 32'b10000000011010000011000101000100; end  // 0,080 -0,997
 944 : begin twid_im = 32'b00001100100010111101001101011110; twid_re = 32'b10000000100111011100100101110010; end  // 0,098 -0,995
 945 : begin twid_im = 32'b00001110111000111000011101100110; twid_re = 32'b10000000110111100110111001001101; end  // 0,116 -0,993
 946 : begin twid_im = 32'b00010001001110011111000011001111; twid_re = 32'b10000001001010100001101000111011; end  // 0,135 -0,991
 947 : begin twid_im = 32'b00010011100011101101101110110001; twid_re = 32'b10000001100000001100011010101010; end  // 0,153 -0,988
 948 : begin twid_im = 32'b00010101111000100001010001000100; twid_re = 32'b10000001111000100110110000010111; end  // 0,171 -0,985
 949 : begin twid_im = 32'b00011000001100110110011011101000; twid_re = 32'b10000010010011110000001000001001; end  // 0,189 -0,982
 950 : begin twid_im = 32'b00011010100000101010000000100101; twid_re = 32'b10000010110001100111111100010101; end  // 0,207 -0,978
 951 : begin twid_im = 32'b00011100110011111000110010110011; twid_re = 32'b10000011010010001101100011011101; end  // 0,225 -0,974
 952 : begin twid_im = 32'b00011111000110011111100101111011; twid_re = 32'b10000011110101100000010000010011; end  // 0,243 -0,970
 953 : begin twid_im = 32'b00100001011000011011001110011111; twid_re = 32'b10000100011011011111010001111000; end  // 0,261 -0,965
 954 : begin twid_im = 32'b00100011101001101000100001111110; twid_re = 32'b10000101000100001001110011011101; end  // 0,279 -0,960
 955 : begin twid_im = 32'b00100101111010000100010110110110; twid_re = 32'b10000101101111011110111100101000; end  // 0,296 -0,955
 956 : begin twid_im = 32'b00101000001001101011100100101000; twid_re = 32'b10000110011101011101110001010000; end  // 0,314 -0,950
 957 : begin twid_im = 32'b00101010011000011011000100000001; twid_re = 32'b10000111001110000101010001011111; end  // 0,331 -0,944
 958 : begin twid_im = 32'b00101100100110001111101110111010; twid_re = 32'b10001000000001010100011001111000; end  // 0,348 -0,937
 959 : begin twid_im = 32'b00101110110011000110100000011110; twid_re = 32'b10001000110111001010000011010100; end  // 0,366 -0,931
 960 : begin twid_im = 32'b00110000111110111100010101001101; twid_re = 32'b10001001101111100101000011000100; end  // 0,383 -0,924
 961 : begin twid_im = 32'b00110011001001101110001011000010; twid_re = 32'b10001010101010100100001010110101; end  // 0,400 -0,917
 962 : begin twid_im = 32'b00110101010011011001000001010110; twid_re = 32'b10001011101000000110001000110000; end  // 0,416 -0,909
 963 : begin twid_im = 32'b00110111011011111001111001000110; twid_re = 32'b10001100101000001001100111011011; end  // 0,433 -0,901
 964 : begin twid_im = 32'b00111001100011001101110100110010; twid_re = 32'b10001101101010101101001101111100; end  // 0,450 -0,893
 965 : begin twid_im = 32'b00111011101001010001111000101001; twid_re = 32'b10001110101111101111011111111100; end  // 0,466 -0,885
 966 : begin twid_im = 32'b00111101101110000011001010100101; twid_re = 32'b10001111110111001110111101100111; end  // 0,482 -0,876
 967 : begin twid_im = 32'b00111111110001011110110010010111; twid_re = 32'b10010001000001001010000011101111; end  // 0,498 -0,867
 968 : begin twid_im = 32'b01000001110011100001111001100100; twid_re = 32'b10010010001101011111001011101100; end  // 0,514 -0,858
 969 : begin twid_im = 32'b01000011110100001001101011101100; twid_re = 32'b10010011011100001100101011100101; end  // 0,530 -0,848
 970 : begin twid_im = 32'b01000101110011010011010110001111; twid_re = 32'b10010100101101010000110110001000; end  // 0,545 -0,838
 971 : begin twid_im = 32'b01000111110000111100001000101110; twid_re = 32'b10010110000000101001111010110110; end  // 0,561 -0,828
 972 : begin twid_im = 32'b01001001101101000001010100110011; twid_re = 32'b10010111010110010110000110000000; end  // 0,576 -0,818
 973 : begin twid_im = 32'b01001011100111100000001110001111; twid_re = 32'b10011000101110010011100000101001; end  // 0,591 -0,807
 974 : begin twid_im = 32'b01001101100000010110001011000011; twid_re = 32'b10011010001000100000010000101110; end  // 0,606 -0,796
 975 : begin twid_im = 32'b01001111010111100000100011100010; twid_re = 32'b10011011100100111010011001000001; end  // 0,620 -0,785
 976 : begin twid_im = 32'b01010001001100111100110010010100; twid_re = 32'b10011101000011011111111001010100; end  // 0,634 -0,773
 977 : begin twid_im = 32'b01010011000000101000010100010111; twid_re = 32'b10011110100100001110101110010101; end  // 0,649 -0,761
 978 : begin twid_im = 32'b01010100110010100000101001001010; twid_re = 32'b10100000000111000100110001110011; end  // 0,662 -0,749
 979 : begin twid_im = 32'b01010110100010100011010010101001; twid_re = 32'b10100001101011111111111010100011; end  // 0,676 -0,737
 980 : begin twid_im = 32'b01011000010000101101110101010100; twid_re = 32'b10100011010010111101111100100001; end  // 0,690 -0,724
 981 : begin twid_im = 32'b01011001111100111101111000010010; twid_re = 32'b10100100111011111100101000110010; end  // 0,703 -0,711
 982 : begin twid_im = 32'b01011011100111010001000101010011; twid_re = 32'b10100110100110111001101101101001; end  // 0,716 -0,698
 983 : begin twid_im = 32'b01011101001111100101001000110110; twid_re = 32'b10101000010011110010110110101011; end  // 0,728 -0,685
 984 : begin twid_im = 32'b01011110110101110111110010001001; twid_re = 32'b10101010000010100101101100101110; end  // 0,741 -0,672
 985 : begin twid_im = 32'b01100000011010000110110011001110; twid_re = 32'b10101011110011001111110110000011; end  // 0,753 -0,658
 986 : begin twid_im = 32'b01100001111100010000000000111110; twid_re = 32'b10101101100101101110110110010010; end  // 0,765 -0,644
 987 : begin twid_im = 32'b01100011011100010001010011001100; twid_re = 32'b10101111011010000000001110100010; end  // 0,777 -0,630
 988 : begin twid_im = 32'b01100100111010001000100100100101; twid_re = 32'b10110001010000000001011101011100; end  // 0,788 -0,615
 989 : begin twid_im = 32'b01100110010101110011110010111011; twid_re = 32'b10110011000111101111111111001100; end  // 0,800 -0,601
 990 : begin twid_im = 32'b01100111101111010000111110111100; twid_re = 32'b10110101000001001001001101101001; end  // 0,810 -0,586
 991 : begin twid_im = 32'b01101001000110011110001100011111; twid_re = 32'b10110110111100001010100000010010; end  // 0,821 -0,571
 992 : begin twid_im = 32'b01101010011011011001100010100011; twid_re = 32'b10111000111000110001001100011010; end  // 0,831 -0,556
 993 : begin twid_im = 32'b01101011101110000001001011010000; twid_re = 32'b10111010110110111010100101000100; end  // 0,842 -0,540
 994 : begin twid_im = 32'b01101100111110010011010011111011; twid_re = 32'b10111100110110100011111011001011; end  // 0,851 -0,525
 995 : begin twid_im = 32'b01101110001100001110001101001001; twid_re = 32'b10111110110111101010011101100110; end  // 0,861 -0,509
 996 : begin twid_im = 32'b01101111010111110000001010110001; twid_re = 32'b11000000111010001011011001001001; end  // 0,870 -0,493
 997 : begin twid_im = 32'b01110000100000110111100011111110; twid_re = 32'b11000010111110000011111000101011; end  // 0,879 -0,477
 998 : begin twid_im = 32'b01110001100111100010110011010001; twid_re = 32'b11000101000011010001000101001001; end  // 0,888 -0,461
 999 : begin twid_im = 32'b01110010101011110000010110100110; twid_re = 32'b11000111001001110000000101101101; end  // 0,896 -0,444
1000 : begin twid_im = 32'b01110011101101011110101111010000; twid_re = 32'b11001001010001011101111111101101; end  // 0,904 -0,428
1001 : begin twid_im = 32'b01110100101100101100100010000011; twid_re = 32'b11001011011010010111110110110001; end  // 0,912 -0,411
1002 : begin twid_im = 32'b01110101101001011000010111001110; twid_re = 32'b11001101100100011010101100111001; end  // 0,919 -0,394
1003 : begin twid_im = 32'b01110110100011100000111010100101; twid_re = 32'b11001111101111100011100010100000; end  // 0,926 -0,377
1004 : begin twid_im = 32'b01110111011011000100111011011010; twid_re = 32'b11010001111011101111010110011110; end  // 0,933 -0,360
1005 : begin twid_im = 32'b01111000010000000011001100101000; twid_re = 32'b11010100001000111011000110010001; end  // 0,939 -0,343
1006 : begin twid_im = 32'b01111001000010011010100100101100; twid_re = 32'b11010110010111000011101101111011; end  // 0,946 -0,325
1007 : begin twid_im = 32'b01111001110010001001111101101101; twid_re = 32'b11011000100110000110001000001100; end  // 0,951 -0,308
1008 : begin twid_im = 32'b01111010011111010000010101011010; twid_re = 32'b11011010110101111111001110100011; end  // 0,957 -0,290
1009 : begin twid_im = 32'b01111011001001101100101101001110; twid_re = 32'b11011101000110101011111001010001; end  // 0,962 -0,273
1010 : begin twid_im = 32'b01111011110001011110001010001111; twid_re = 32'b11011111011000001000111111100100; end  // 0,967 -0,255
1011 : begin twid_im = 32'b01111100010110100011110101001111; twid_re = 32'b11100001101010010011010111100010; end  // 0,972 -0,237
1012 : begin twid_im = 32'b01111100111000111100111010110001; twid_re = 32'b11100011111101000111110110010110; end  // 0,976 -0,219
1013 : begin twid_im = 32'b01111101011000101000101011000101; twid_re = 32'b11100110010000100011010000001101; end  // 0,980 -0,201
1014 : begin twid_im = 32'b01111101110101100110011010001110; twid_re = 32'b11101000100100100010011000100010; end  // 0,983 -0,183
1015 : begin twid_im = 32'b01111110001111110101011111111110; twid_re = 32'b11101010111001000010000001111011; end  // 0,986 -0,165
1016 : begin twid_im = 32'b01111110100111010101010111111011; twid_re = 32'b11101101001101111110111110010010; end  // 0,989 -0,147
1017 : begin twid_im = 32'b01111110111100000101100001011111; twid_re = 32'b11101111100011010101111110111000; end  // 0,992 -0,128
1018 : begin twid_im = 32'b01111111001110000101011111110101; twid_re = 32'b11110001111001000011110100011100; end  // 0,994 -0,110
1019 : begin twid_im = 32'b01111111011101010100111001111111; twid_re = 32'b11110100001111000101001111001011; end  // 0,996 -0,092
1020 : begin twid_im = 32'b01111111101001110011011010110011; twid_re = 32'b11110110100101010110111110110111; end  // 0,997 -0,074
1021 : begin twid_im = 32'b01111111110011100000110000111101; twid_re = 32'b11111000111011110101110010111011; end  // 0,998 -0,055
1022 : begin twid_im = 32'b01111111111010011100101110111111; twid_re = 32'b11111011010010011110011010100011; end  // 0,999 -0,037
1023 : begin twid_im = 32'b01111111111110100111001011010000; twid_re = 32'b11111101101001001101100100101001; end  // 1,000 -0,018
    endcase 
endmodule 


`timescale 1ns/10ps

module COREFFT_C0_COREFFT_C0_0_twidLut_stage_4 (index, twid_im, twid_re);
  input[7:0] index;
  output [31:0] twid_im, twid_re;
  reg    signed [31:0] twid_im, twid_re;

  always @ (index) 
    case (index) 
   0 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   1 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   2 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   3 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   4 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   5 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   6 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   7 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   8 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   9 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  10 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  11 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  12 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  13 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  14 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  15 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  16 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  17 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  18 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  19 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  20 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  21 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  22 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  23 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  24 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  25 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  26 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  27 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  28 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  29 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  30 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  31 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  32 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  33 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  34 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  35 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  36 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  37 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  38 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  39 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  40 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  41 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  42 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  43 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  44 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  45 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  46 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  47 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  48 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  49 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  50 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  51 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  52 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  53 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  54 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  55 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  56 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  57 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  58 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  59 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  60 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  61 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  62 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  63 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  64 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  65 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b01111111110110001000011110001101; end  //-0,049  0,999
  66 : begin twid_im = 32'b11110011011101000010110010100010; twid_re = 32'b01111111011000100011011010001110; end  //-0,098  0,995
  67 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b01111110100111010101010111111011; end  //-0,147  0,989
  68 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b01111101100010100101111100111111; end  //-0,195  0,981
  69 : begin twid_im = 32'b11100000111001100000011010000101; twid_re = 32'b01111100001010011111101111101101; end  //-0,243  0,970
  70 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
  71 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b01111000100001001000010000010011; end  //-0,337  0,942
  72 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b01110110010000011010111100111100; end  //-0,383  0,924
  73 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b01110011101101011110101111010000; end  //-0,428  0,904
  74 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b01110000111000101100101111000101; end  //-0,471  0,882
  75 : begin twid_im = 32'b10111110001100011110000110011100; twid_re = 32'b01101101110010100000110100010100; end  //-0,514  0,858
  76 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
  77 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b01100110110011111000000100011111; end  //-0,596  0,803
  78 : begin twid_im = 32'b10101110110011000011001101101100; twid_re = 32'b01100010111100100000000110101100; end  //-0,634  0,773
  79 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b01011110110101110111110010001001; end  //-0,672  0,741
  80 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
  81 : begin twid_im = 32'b10100001001010001000001101110111; twid_re = 32'b01010101111101011010010011010010; end  //-0,741  0,672
  82 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
  83 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b01001100001111111101111111110011; end  //-0,803  0,596
  84 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b01000111000111001110110011100110; end  //-0,831  0,556
  85 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b01000001110011100001111001100100; end  //-0,858  0,514
  86 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b00111100010101101011101001110000; end  //-0,882  0,471
  87 : begin twid_im = 32'b10001100010010100001010000110000; twid_re = 32'b00110110101110100010000000010011; end  //-0,904  0,428
  88 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
  89 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b00101011000111110011010011101011; end  //-0,942  0,337
  90 : begin twid_im = 32'b10000101100000101111101010100110; twid_re = 32'b00100101001010000000110001011101; end  //-0,957  0,290
  91 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b00011111000110011111100101111011; end  //-0,970  0,243
  92 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b00011000111110001011100000111100; end  //-0,981  0,195
  93 : begin twid_im = 32'b10000001011000101010101000000101; twid_re = 32'b00010010110010000001000001101110; end  //-0,989  0,147
  94 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
  95 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b00000110010001111101100101111100; end  //-0,999  0,049
  96 : begin twid_im = 32'b10000000000000000000000000000001; twid_re = 32'b00000000000000000000000000000000; end  //-1,000  0,000
  97 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b11111001101110000010011010000100; end  //-0,999 -0,049
  98 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b11110011011101000010110010100010; end  //-0,995 -0,098
  99 : begin twid_im = 32'b10000001011000101010101000000101; twid_re = 32'b11101101001101111110111110010010; end  //-0,989 -0,147
 100 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b11100111000001110100011111000100; end  //-0,981 -0,195
 101 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b11100000111001100000011010000101; end  //-0,970 -0,243
 102 : begin twid_im = 32'b10000101100000101111101010100110; twid_re = 32'b11011010110101111111001110100011; end  //-0,957 -0,290
 103 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b11010100111000001100101100010101; end  //-0,942 -0,337
 104 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b11001111000001000011101010110011; end  //-0,924 -0,383
 105 : begin twid_im = 32'b10001100010010100001010000110000; twid_re = 32'b11001001010001011101111111101101; end  //-0,904 -0,428
 106 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b11000011101010010100010110010000; end  //-0,882 -0,471
 107 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b10111110001100011110000110011100; end  //-0,858 -0,514
 108 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b10111000111000110001001100011010; end  //-0,831 -0,556
 109 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b10110011110000000010000000001101; end  //-0,803 -0,596
 110 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b10101110110011000011001101101100; end  //-0,773 -0,634
 111 : begin twid_im = 32'b10100001001010001000001101110111; twid_re = 32'b10101010000010100101101100101110; end  //-0,741 -0,672
 112 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
 113 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b10100001001010001000001101110111; end  //-0,672 -0,741
 114 : begin twid_im = 32'b10101110110011000011001101101100; twid_re = 32'b10011101000011011111111001010100; end  //-0,634 -0,773
 115 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b10011001001100000111111011100001; end  //-0,596 -0,803
 116 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b10010101100100100110011101011101; end  //-0,556 -0,831
 117 : begin twid_im = 32'b10111110001100011110000110011100; twid_re = 32'b10010010001101011111001011101100; end  //-0,514 -0,858
 118 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b10001111000111010011010000111011; end  //-0,471 -0,882
 119 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b10001100010010100001010000110000; end  //-0,428 -0,904
 120 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b10001001101111100101000011000100; end  //-0,383 -0,924
 121 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b10000111011110110111101111101101; end  //-0,337 -0,942
 122 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b10000101100000101111101010100110; end  //-0,290 -0,957
 123 : begin twid_im = 32'b11100000111001100000011010000101; twid_re = 32'b10000011110101100000010000010011; end  //-0,243 -0,970
 124 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b10000010011101011010000011000001; end  //-0,195 -0,981
 125 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b10000001011000101010101000000101; end  //-0,147 -0,989
 126 : begin twid_im = 32'b11110011011101000010110010100010; twid_re = 32'b10000000100111011100100101110010; end  //-0,098 -0,995
 127 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b10000000001001110111100001110011; end  //-0,049 -0,999
 128 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 129 : begin twid_im = 32'b11111100110110111101010101000001; twid_re = 32'b01111111111101100010000110000001; end  //-0,025  1,000
 130 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b01111111110110001000011110001101; end  //-0,049  0,999
 131 : begin twid_im = 32'b11110110100101010110111110110111; twid_re = 32'b01111111101001110011011010110011; end  //-0,074  0,997
 132 : begin twid_im = 32'b11110011011101000010110010100010; twid_re = 32'b01111111011000100011011010001110; end  //-0,098  0,995
 133 : begin twid_im = 32'b11110000010101001101100011010101; twid_re = 32'b01111111000010011001000111000011; end  //-0,122  0,992
 134 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b01111110100111010101010111111011; end  //-0,147  0,989
 135 : begin twid_im = 32'b11101010000111011110101110111100; twid_re = 32'b01111110000111011001001111101001; end  //-0,171  0,985
 136 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b01111101100010100101111100111111; end  //-0,195  0,981
 137 : begin twid_im = 32'b11100011111101000111110110010110; twid_re = 32'b01111100111000111100111010110001; end  //-0,219  0,976
 138 : begin twid_im = 32'b11100000111001100000011010000101; twid_re = 32'b01111100001010011111101111101101; end  //-0,243  0,970
 139 : begin twid_im = 32'b11011101110111000101101100111011; twid_re = 32'b01111011010111010000001110011101; end  //-0,267  0,964
 140 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
 141 : begin twid_im = 32'b11010111110110010100011011011000; twid_re = 32'b01111001100010100010001110110000; end  //-0,314  0,950
 142 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b01111000100001001000010000010011; end  //-0,337  0,942
 143 : begin twid_im = 32'b11010001111011101111010110011110; twid_re = 32'b01110111011011000100111011011010; end  //-0,360  0,933
 144 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b01110110010000011010111100111100; end  //-0,383  0,924
 145 : begin twid_im = 32'b11001100001000010000110101111001; twid_re = 32'b01110101000001001101001101000100; end  //-0,405  0,914
 146 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b01110011101101011110101111010000; end  //-0,428  0,904
 147 : begin twid_im = 32'b11000110011100110010001011001110; twid_re = 32'b01110010010101010010110010000100; end  //-0,450  0,893
 148 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b01110000111000101100101111000101; end  //-0,471  0,882
 149 : begin twid_im = 32'b11000000111010001011011001001001; twid_re = 32'b01101111010111110000001010110001; end  //-0,493  0,870
 150 : begin twid_im = 32'b10111110001100011110000110011100; twid_re = 32'b01101101110010100000110100010100; end  //-0,514  0,858
 151 : begin twid_im = 32'b10111011100001010011001010110000; twid_re = 32'b01101100001001000010100101011111; end  //-0,535  0,845
 152 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
 153 : begin twid_im = 32'b10110110010010111110101011001101; twid_re = 32'b01101000101001101001111010000000; end  //-0,576  0,818
 154 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b01100110110011111000000100011111; end  //-0,596  0,803
 155 : begin twid_im = 32'b10110001010000000001011101011100; twid_re = 32'b01100100111010001000100100100101; end  //-0,615  0,788
 156 : begin twid_im = 32'b10101110110011000011001101101100; twid_re = 32'b01100010111100100000000110101100; end  //-0,634  0,773
 157 : begin twid_im = 32'b10101100011001001101010100010001; twid_re = 32'b01100000111011000011100000101111; end  //-0,653  0,757
 158 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b01011110110101110111110010001001; end  //-0,672  0,741
 159 : begin twid_im = 32'b10100111101111010010001010101100; twid_re = 32'b01011100101101000010000011011111; end  //-0,690  0,724
 160 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
 161 : begin twid_im = 32'b10100011010010111101111100100001; twid_re = 32'b01011000010000101101110101010100; end  //-0,724  0,690
 162 : begin twid_im = 32'b10100001001010001000001101110111; twid_re = 32'b01010101111101011010010011010010; end  //-0,741  0,672
 163 : begin twid_im = 32'b10011111000100111100011111010001; twid_re = 32'b01010011100110110010101011101111; end  //-0,757  0,653
 164 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
 165 : begin twid_im = 32'b10011011000101110111011011011011; twid_re = 32'b01001110101111111110100010100100; end  //-0,788  0,615
 166 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b01001100001111111101111111110011; end  //-0,803  0,596
 167 : begin twid_im = 32'b10010111010110010110000110000000; twid_re = 32'b01001001101101000001010100110011; end  //-0,818  0,576
 168 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b01000111000111001110110011100110; end  //-0,831  0,556
 169 : begin twid_im = 32'b10010011110110111101011010100001; twid_re = 32'b01000100011110101100110101010000; end  //-0,845  0,535
 170 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b01000001110011100001111001100100; end  //-0,858  0,514
 171 : begin twid_im = 32'b10010000101000001111110101001111; twid_re = 32'b00111111000101110100100110110111; end  //-0,870  0,493
 172 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b00111100010101101011101001110000; end  //-0,882  0,471
 173 : begin twid_im = 32'b10001101101010101101001101111100; twid_re = 32'b00111001100011001101110100110010; end  //-0,893  0,450
 174 : begin twid_im = 32'b10001100010010100001010000110000; twid_re = 32'b00110110101110100010000000010011; end  //-0,904  0,428
 175 : begin twid_im = 32'b10001010111110110010110010111100; twid_re = 32'b00110011110111101111001010000111; end  //-0,914  0,405
 176 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
 177 : begin twid_im = 32'b10001000100100111011000100100110; twid_re = 32'b00101110000100010000101001100010; end  //-0,933  0,360
 178 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b00101011000111110011010011101011; end  //-0,942  0,337
 179 : begin twid_im = 32'b10000110011101011101110001010000; twid_re = 32'b00101000001001101011100100101000; end  //-0,950  0,314
 180 : begin twid_im = 32'b10000101100000101111101010100110; twid_re = 32'b00100101001010000000110001011101; end  //-0,957  0,290
 181 : begin twid_im = 32'b10000100101000101111110001100011; twid_re = 32'b00100010001000111010010011000101; end  //-0,964  0,267
 182 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b00011111000110011111100101111011; end  //-0,970  0,243
 183 : begin twid_im = 32'b10000011000111000011000101001111; twid_re = 32'b00011100000010111000001001101010; end  //-0,976  0,219
 184 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b00011000111110001011100000111100; end  //-0,981  0,195
 185 : begin twid_im = 32'b10000001111000100110110000010111; twid_re = 32'b00010101111000100001010001000100; end  //-0,985  0,171
 186 : begin twid_im = 32'b10000001011000101010101000000101; twid_re = 32'b00010010110010000001000001101110; end  //-0,989  0,147
 187 : begin twid_im = 32'b10000000111101100110111000111101; twid_re = 32'b00001111101010110010011100101011; end  //-0,992  0,122
 188 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
 189 : begin twid_im = 32'b10000000010110001100100101001101; twid_re = 32'b00001001011010101001000001001001; end  //-0,997  0,074
 190 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b00000110010001111101100101111100; end  //-0,999  0,049
 191 : begin twid_im = 32'b10000000000010011101111001111111; twid_re = 32'b00000011001001000010101010111111; end  //-1,000  0,025
 192 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
 193 : begin twid_im = 32'b11110110100101010110111110110111; twid_re = 32'b01111111101001110011011010110011; end  //-0,074  0,997
 194 : begin twid_im = 32'b11101101001101111110111110010010; twid_re = 32'b01111110100111010101010111111011; end  //-0,147  0,989
 195 : begin twid_im = 32'b11100011111101000111110110010110; twid_re = 32'b01111100111000111100111010110001; end  //-0,219  0,976
 196 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
 197 : begin twid_im = 32'b11010001111011101111010110011110; twid_re = 32'b01110111011011000100111011011010; end  //-0,360  0,933
 198 : begin twid_im = 32'b11001001010001011101111111101101; twid_re = 32'b01110011101101011110101111010000; end  //-0,428  0,904
 199 : begin twid_im = 32'b11000000111010001011011001001001; twid_re = 32'b01101111010111110000001010110001; end  //-0,493  0,870
 200 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
 201 : begin twid_im = 32'b10110001010000000001011101011100; twid_re = 32'b01100100111010001000100100100101; end  //-0,615  0,788
 202 : begin twid_im = 32'b10101010000010100101101100101110; twid_re = 32'b01011110110101110111110010001001; end  //-0,672  0,741
 203 : begin twid_im = 32'b10100011010010111101111100100001; twid_re = 32'b01011000010000101101110101010100; end  //-0,724  0,690
 204 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
 205 : begin twid_im = 32'b10010111010110010110000110000000; twid_re = 32'b01001001101101000001010100110011; end  //-0,818  0,576
 206 : begin twid_im = 32'b10010010001101011111001011101100; twid_re = 32'b01000001110011100001111001100100; end  //-0,858  0,514
 207 : begin twid_im = 32'b10001101101010101101001101111100; twid_re = 32'b00111001100011001101110100110010; end  //-0,893  0,450
 208 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
 209 : begin twid_im = 32'b10000110011101011101110001010000; twid_re = 32'b00101000001001101011100100101000; end  //-0,950  0,314
 210 : begin twid_im = 32'b10000011110101100000010000010011; twid_re = 32'b00011111000110011111100101111011; end  //-0,970  0,243
 211 : begin twid_im = 32'b10000001111000100110110000010111; twid_re = 32'b00010101111000100001010001000100; end  //-0,985  0,171
 212 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
 213 : begin twid_im = 32'b10000000000010011101111001111111; twid_re = 32'b00000011001001000010101010111111; end  //-1,000  0,025
 214 : begin twid_im = 32'b10000000001001110111100001110011; twid_re = 32'b11111001101110000010011010000100; end  //-0,999 -0,049
 215 : begin twid_im = 32'b10000000111101100110111000111101; twid_re = 32'b11110000010101001101100011010101; end  //-0,992 -0,122
 216 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b11100111000001110100011111000100; end  //-0,981 -0,195
 217 : begin twid_im = 32'b10000100101000101111110001100011; twid_re = 32'b11011101110111000101101100111011; end  //-0,964 -0,267
 218 : begin twid_im = 32'b10000111011110110111101111101101; twid_re = 32'b11010100111000001100101100010101; end  //-0,942 -0,337
 219 : begin twid_im = 32'b10001010111110110010110010111100; twid_re = 32'b11001100001000010000110101111001; end  //-0,914 -0,405
 220 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b11000011101010010100010110010000; end  //-0,882 -0,471
 221 : begin twid_im = 32'b10010011110110111101011010100001; twid_re = 32'b10111011100001010011001010110000; end  //-0,845 -0,535
 222 : begin twid_im = 32'b10011001001100000111111011100001; twid_re = 32'b10110011110000000010000000001101; end  //-0,803 -0,596
 223 : begin twid_im = 32'b10011111000100111100011111010001; twid_re = 32'b10101100011001001101010100010001; end  //-0,757 -0,653
 224 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
 225 : begin twid_im = 32'b10101100011001001101010100010001; twid_re = 32'b10011111000100111100011111010001; end  //-0,653 -0,757
 226 : begin twid_im = 32'b10110011110000000010000000001101; twid_re = 32'b10011001001100000111111011100001; end  //-0,596 -0,803
 227 : begin twid_im = 32'b10111011100001010011001010110000; twid_re = 32'b10010011110110111101011010100001; end  //-0,535 -0,845
 228 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b10001111000111010011010000111011; end  //-0,471 -0,882
 229 : begin twid_im = 32'b11001100001000010000110101111001; twid_re = 32'b10001010111110110010110010111100; end  //-0,405 -0,914
 230 : begin twid_im = 32'b11010100111000001100101100010101; twid_re = 32'b10000111011110110111101111101101; end  //-0,337 -0,942
 231 : begin twid_im = 32'b11011101110111000101101100111011; twid_re = 32'b10000100101000101111110001100011; end  //-0,267 -0,964
 232 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b10000010011101011010000011000001; end  //-0,195 -0,981
 233 : begin twid_im = 32'b11110000010101001101100011010101; twid_re = 32'b10000000111101100110111000111101; end  //-0,122 -0,992
 234 : begin twid_im = 32'b11111001101110000010011010000100; twid_re = 32'b10000000001001110111100001110011; end  //-0,049 -0,999
 235 : begin twid_im = 32'b00000011001001000010101010111111; twid_re = 32'b10000000000010011101111001111111; end  // 0,025 -1,000
 236 : begin twid_im = 32'b00001100100010111101001101011110; twid_re = 32'b10000000100111011100100101110010; end  // 0,098 -0,995
 237 : begin twid_im = 32'b00010101111000100001010001000100; twid_re = 32'b10000001111000100110110000010111; end  // 0,171 -0,985
 238 : begin twid_im = 32'b00011111000110011111100101111011; twid_re = 32'b10000011110101100000010000010011; end  // 0,243 -0,970
 239 : begin twid_im = 32'b00101000001001101011100100101000; twid_re = 32'b10000110011101011101110001010000; end  // 0,314 -0,950
 240 : begin twid_im = 32'b00110000111110111100010101001101; twid_re = 32'b10001001101111100101000011000100; end  // 0,383 -0,924
 241 : begin twid_im = 32'b00111001100011001101110100110010; twid_re = 32'b10001101101010101101001101111100; end  // 0,450 -0,893
 242 : begin twid_im = 32'b01000001110011100001111001100100; twid_re = 32'b10010010001101011111001011101100; end  // 0,514 -0,858
 243 : begin twid_im = 32'b01001001101101000001010100110011; twid_re = 32'b10010111010110010110000110000000; end  // 0,576 -0,818
 244 : begin twid_im = 32'b01010001001100111100110010010100; twid_re = 32'b10011101000011011111111001010100; end  // 0,634 -0,773
 245 : begin twid_im = 32'b01011000010000101101110101010100; twid_re = 32'b10100011010010111101111100100001; end  // 0,690 -0,724
 246 : begin twid_im = 32'b01011110110101110111110010001001; twid_re = 32'b10101010000010100101101100101110; end  // 0,741 -0,672
 247 : begin twid_im = 32'b01100100111010001000100100100101; twid_re = 32'b10110001010000000001011101011100; end  // 0,788 -0,615
 248 : begin twid_im = 32'b01101010011011011001100010100011; twid_re = 32'b10111000111000110001001100011010; end  // 0,831 -0,556
 249 : begin twid_im = 32'b01101111010111110000001010110001; twid_re = 32'b11000000111010001011011001001001; end  // 0,870 -0,493
 250 : begin twid_im = 32'b01110011101101011110101111010000; twid_re = 32'b11001001010001011101111111101101; end  // 0,904 -0,428
 251 : begin twid_im = 32'b01110111011011000100111011011010; twid_re = 32'b11010001111011101111010110011110; end  // 0,933 -0,360
 252 : begin twid_im = 32'b01111010011111010000010101011010; twid_re = 32'b11011010110101111111001110100011; end  // 0,957 -0,290
 253 : begin twid_im = 32'b01111100111000111100111010110001; twid_re = 32'b11100011111101000111110110010110; end  // 0,976 -0,219
 254 : begin twid_im = 32'b01111110100111010101010111111011; twid_re = 32'b11101101001101111110111110010010; end  // 0,989 -0,147
 255 : begin twid_im = 32'b01111111101001110011011010110011; twid_re = 32'b11110110100101010110111110110111; end  // 0,997 -0,074
    endcase 
endmodule 


`timescale 1ns/10ps

module COREFFT_C0_COREFFT_C0_0_twidLut_stage_6 (index, twid_im, twid_re);
  input[5:0] index;
  output [31:0] twid_im, twid_re;
  reg    signed [31:0] twid_im, twid_re;

  always @ (index) 
    case (index) 
   0 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   1 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   2 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   3 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   4 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   5 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   6 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   7 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   8 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   9 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  10 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  11 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  12 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  13 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  14 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  15 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  16 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  17 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b01111101100010100101111100111111; end  //-0,195  0,981
  18 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b01110110010000011010111100111100; end  //-0,383  0,924
  19 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
  20 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
  21 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b01000111000111001110110011100110; end  //-0,831  0,556
  22 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
  23 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b00011000111110001011100000111100; end  //-0,981  0,195
  24 : begin twid_im = 32'b10000000000000000000000000000001; twid_re = 32'b00000000000000000000000000000000; end  //-1,000  0,000
  25 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b11100111000001110100011111000100; end  //-0,981 -0,195
  26 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b11001111000001000011101010110011; end  //-0,924 -0,383
  27 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b10111000111000110001001100011010; end  //-0,831 -0,556
  28 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
  29 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b10010101100100100110011101011101; end  //-0,556 -0,831
  30 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b10001001101111100101000011000100; end  //-0,383 -0,924
  31 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b10000010011101011010000011000001; end  //-0,195 -0,981
  32 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  33 : begin twid_im = 32'b11110011011101000010110010100010; twid_re = 32'b01111111011000100011011010001110; end  //-0,098  0,995
  34 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b01111101100010100101111100111111; end  //-0,195  0,981
  35 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
  36 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b01110110010000011010111100111100; end  //-0,383  0,924
  37 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b01110000111000101100101111000101; end  //-0,471  0,882
  38 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
  39 : begin twid_im = 32'b10101110110011000011001101101100; twid_re = 32'b01100010111100100000000110101100; end  //-0,634  0,773
  40 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
  41 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
  42 : begin twid_im = 32'b10010101100100100110011101011101; twid_re = 32'b01000111000111001110110011100110; end  //-0,831  0,556
  43 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b00111100010101101011101001110000; end  //-0,882  0,471
  44 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
  45 : begin twid_im = 32'b10000101100000101111101010100110; twid_re = 32'b00100101001010000000110001011101; end  //-0,957  0,290
  46 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b00011000111110001011100000111100; end  //-0,981  0,195
  47 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
  48 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  49 : begin twid_im = 32'b11011010110101111111001110100011; twid_re = 32'b01111010011111010000010101011010; end  //-0,290  0,957
  50 : begin twid_im = 32'b10111000111000110001001100011010; twid_re = 32'b01101010011011011001100010100011; end  //-0,556  0,831
  51 : begin twid_im = 32'b10011101000011011111111001010100; twid_re = 32'b01010001001100111100110010010100; end  //-0,773  0,634
  52 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
  53 : begin twid_im = 32'b10000000100111011100100101110010; twid_re = 32'b00001100100010111101001101011110; end  //-0,995  0,098
  54 : begin twid_im = 32'b10000010011101011010000011000001; twid_re = 32'b11100111000001110100011111000100; end  //-0,981 -0,195
  55 : begin twid_im = 32'b10001111000111010011010000111011; twid_re = 32'b11000011101010010100010110010000; end  //-0,882 -0,471
  56 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
  57 : begin twid_im = 32'b11000011101010010100010110010000; twid_re = 32'b10001111000111010011010000111011; end  //-0,471 -0,882
  58 : begin twid_im = 32'b11100111000001110100011111000100; twid_re = 32'b10000010011101011010000011000001; end  //-0,195 -0,981
  59 : begin twid_im = 32'b00001100100010111101001101011110; twid_re = 32'b10000000100111011100100101110010; end  // 0,098 -0,995
  60 : begin twid_im = 32'b00110000111110111100010101001101; twid_re = 32'b10001001101111100101000011000100; end  // 0,383 -0,924
  61 : begin twid_im = 32'b01010001001100111100110010010100; twid_re = 32'b10011101000011011111111001010100; end  // 0,634 -0,773
  62 : begin twid_im = 32'b01101010011011011001100010100011; twid_re = 32'b10111000111000110001001100011010; end  // 0,831 -0,556
  63 : begin twid_im = 32'b01111010011111010000010101011010; twid_re = 32'b11011010110101111111001110100011; end  // 0,957 -0,290
    endcase 
endmodule 


`timescale 1ns/10ps

module COREFFT_C0_COREFFT_C0_0_twidLut_stage_8 (index, twid_im, twid_re);
  input[3:0] index;
  output [31:0] twid_im, twid_re;
  reg    signed [31:0] twid_im, twid_re;

  always @ (index) 
    case (index) 
   0 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   1 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   2 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   3 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   4 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   5 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
   6 : begin twid_im = 32'b10000000000000000000000000000001; twid_re = 32'b00000000000000000000000000000000; end  //-1,000  0,000
   7 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
   8 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
   9 : begin twid_im = 32'b11001111000001000011101010110011; twid_re = 32'b01110110010000011010111100111100; end  //-0,383  0,924
  10 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b01011010100000100111100110011001; end  //-0,707  0,707
  11 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
  12 : begin twid_im = 32'b00000000000000000000000000000000; twid_re = 32'b01111111111111111111111111111111; end  //-0,000  1,000
  13 : begin twid_im = 32'b10001001101111100101000011000100; twid_re = 32'b00110000111110111100010101001101; end  //-0,924  0,383
  14 : begin twid_im = 32'b10100101011111011000011001100111; twid_re = 32'b10100101011111011000011001100111; end  //-0,707 -0,707
  15 : begin twid_im = 32'b00110000111110111100010101001101; twid_re = 32'b10001001101111100101000011000100; end  // 0,383 -0,924
    endcase 
endmodule 


