// -----------------------------------------------------------------------------
//Actel Corporation Proprietary and Confidential
//Copyright 2008 Actel Corporation. All rights reserved.
//
//ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
//ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
//IN ADVANCE IN WRITING.
//
//Description:  CoreFFT RTL 
//              Customized Twiddle Coefficients 
//
//Revision Information:
//Date         Description
//05Nov2009    Initial Release 
//
//SVN Revision Information:
//SVN $Revision: $
//SVN $Data: $
//
//Resolved SARs
//SAR     Date    Who         Description
//
//Notes:

`timescale 1 ns/100 ps

module COREFFT_C0_COREFFT_C0_0_twiddle (A,T);
  parameter TDWIDTH = 16;
  parameter LOGPTS  = 5;

  input	[LOGPTS-2:0]	A;	// Address
  output reg [TDWIDTH-1:0]	T;	// Table output

  always @ (A)
    case (A) // synopsys parallel_case
      9'h0: T=64'b0000000000000000000000000000000001111111111111111111111111111111;  //     0 2147483647
      9'h1: T=64'b1111111100110110111100000111100001111111111111110110001000010101;  // -13176712 2147443221
      9'h2: T=64'b1111111001101101111000101110000001111111111111011000100001011001;  // -26352928 2147321945
      9'h3: T=64'b1111110110100100110110010010100101111111111110100111001011010000;  // -39528151 2147119824
      9'h4: T=64'b1111110011011011110101010100000101111111111101100010000110000001;  // -52701887 2146836865
      9'h5: T=64'b1111110000010010110110010001101001111111111100001001010001110111;  // -65873638 2146473079
      9'h6: T=64'b1111101101001001111001101010001101111111111010011100101110111111;  // -79042909 2146028479
      9'h7: T=64'b1111101010000000111111111100101101111111111000011100011101101010;  // -92209205 2145503082
      9'h8: T=64'b1111100110111000001001101000010001111111110110001000011110001101;  // -105372028 2144896909
      9'h9: T=64'b1111100011101111010111001011101101111111110011100000110000111101;  // -118530885 2144209981
      9'ha: T=64'b1111100000100110101001000110001001111111110000100101010110010101;  // -131685278 2143442325
      9'hb: T=64'b1111011101011101111111110110011001111111101101010110001110110010;  // -144834714 2142593970
      9'hc: T=64'b1111011010010101011011111011011101111111101001110011011010110011;  // -157978697 2141664947
      9'hd: T=64'b1111010111001100111101110100010001111111100101111100111010111100;  // -171116732 2140655292
      9'he: T=64'b1111010100000100100101111111101101111111100001110010101111110010;  // -184248325 2139565042
      9'hf: T=64'b1111010000111100010100111100101101111111011101010100111001111111;  // -197372981 2138394239
      9'h10: T=64'b1111001101110100001011001010001001111111011000100011011010001110;  // -210490206 2137142926
      9'h11: T=64'b1111001010101100001001000110111001111111010011011110010001010000;  // -223599506 2135811152
      9'h12: T=64'b1111000111100100001111010001110001111111001110000101011111110101;  // -236700388 2134398965
      9'h13: T=64'b1111000100011100011110001001101001111111001000011001000110110011;  // -249792358 2132906419
      9'h14: T=64'b1111000001010100110110001101010101111111000010011001000111000011;  // -262874923 2131333571
      9'h15: T=64'b1110111110001101010111111011100001111110111100000101100001011111;  // -275947592 2129680479
      9'h16: T=64'b1110111011000110000011110011000101111110110101011110010111000101;  // -289009871 2127947205
      9'h17: T=64'b1110110111111110111010010010101101111110101110100011101000111000;  // -302061269 2126133816
      9'h18: T=64'b1110110100110111111011111001001001111110100111010101010111111011;  // -315101294 2124240379
      9'h19: T=64'b1110110001110001001001000100111101111110011111110011100101010110;  // -328129457 2122266966
      9'h1a: T=64'b1110101110101010100010010100111101111110010111111110010010010010;  // -341145265 2120213650
      9'h1b: T=64'b1110101011100100001000000111101101111110001111110101011111111110;  // -354148229 2118080510
      9'h1c: T=64'b1110101000011101111010111011110001111110000111011001001111101001;  // -367137860 2115867625
      9'h1d: T=64'b1110100101010111111011001111101101111101111110101001100010100111;  // -380113669 2113575079
      9'h1e: T=64'b1110100010010010001001100010001001111101110101100110011010001110;  // -393075166 2111202958
      9'h1f: T=64'b1110011111001100100110010001100001111101101100001111110111110111;  // -406021864 2108751351
      9'h20: T=64'b1110011100000111010001111100010001111101100010100101111100111111;  // -418953276 2106220351
      9'h21: T=64'b1110011001000010001101000000110101111101011000101000101011000101;  // -431868915 2103610053
      9'h22: T=64'b1110010101111101010111111101101101111101001110011000000011101011;  // -444768293 2100920555
      9'h23: T=64'b1110010010111000110011010001000101111101000011110100001000010111;  // -457650927 2098151959
      9'h24: T=64'b1110001111110100011111011001011001111100111000111100111010110001;  // -470516330 2095304369
      9'h25: T=64'b1110001100110000011100110100110101111100101101110010011100100011;  // -483364019 2092377891
      9'h26: T=64'b1110001001101100101100000001101101111100100010010100101111011101;  // -496193509 2089372637
      9'h27: T=64'b1110000110101001001101011110001001111100010110100011110101001111;  // -509004318 2086288719
      9'h28: T=64'b1110000011100110000001101000010101111100001010011111101111101101;  // -521795963 2083126253
      9'h29: T=64'b1110000000100011001000111110010101111011111110001000100000101111;  // -534567963 2079885359
      9'h2a: T=64'b1101111101100000100011111110010001111011110001011110001010001111;  // -547319836 2076566159
      9'h2b: T=64'b1101111010011110010011000110000101111011100100100000101110001000;  // -560051103 2073168776
      9'h2c: T=64'b1101110111011100010110110011101101111011010111010000001110011101;  // -572761285 2069693341
      9'h2d: T=64'b1101110100011010101111100101000101111011001001101100101101001110;  // -585449903 2066139982
      9'h2e: T=64'b1101110001011001011101111000001001111010111011110110001100100011;  // -598116478 2062508835
      9'h2f: T=64'b1101101110011000100010001010100101111010101101101100101110100011;  // -610760535 2058800035
      9'h30: T=64'b1101101011010111111100111010001101111010011111010000010101011010;  // -623381597 2055013722
      9'h31: T=64'b1101101000010111101110100100101001111010010000100001000011011000;  // -635979190 2051150040
      9'h32: T=64'b1101100101010111110111100111101101111010000001011110111010101100;  // -648552837 2047209132
      9'h33: T=64'b1101100010011000011000100000110001111001110010001001111101101101;  // -661102068 2043191149
      9'h34: T=64'b1101011111011001010001101101100001111001100010100010001110110000;  // -673626408 2039096240
      9'h35: T=64'b1101011100011010100011101011011001111001010010100111110000010001;  // -686125386 2034924561
      9'h36: T=64'b1101011001011100001110110111101101111001000010011010100100101100;  // -698598533 2030676268
      9'h37: T=64'b1101010110011110010011101111111101111000110001111010101110100001;  // -711045377 2026351521
      9'h38: T=64'b1101010011100000110010110001010101111000100001001000010000010011;  // -723465451 2021950483
      9'h39: T=64'b1101010000100011101100011001000101111000010000000011001100101000;  // -735858287 2017473320
      9'h3a: T=64'b1101001101100111000001000100011001110111111110101011100110001000;  // -748223418 2012920200
      9'h3b: T=64'b1101001010101010110001010000010101110111101101000001011111011111;  // -760560379 2008291295
      9'h3c: T=64'b1101000111101110111101011001111001110111011011000100111011011010;  // -772868706 2003586778
      9'h3d: T=64'b1101000100110011100101111110001001110111001000110101111100101100;  // -785147934 1998806828
      9'h3e: T=64'b1101000001111000101011011001111001110110110110010100100110001000;  // -797397602 1993951624
      9'h3f: T=64'b1100111110111110001110001010000001110110100011100000111010100101;  // -809617248 1989021349
      9'h40: T=64'b1100111100000100001110101011001101110110010000011010111100111100;  // -821806413 1984016188
      9'h41: T=64'b1100111001001010101101011010001101110101111101000010110000001010;  // -833964637 1978936330
      9'h42: T=64'b1100110110010001101010110011100101110101101001011000010111001110;  // -846091463 1973781966
      9'h43: T=64'b1100110011011001000111010011111001110101010101011011110101001011;  // -858186434 1968553291
      9'h44: T=64'b1100110000100001000011010111100101110101000001001101001101000100;  // -870249095 1963250500
      9'h45: T=64'b1100101101101001011111011011000101110100101100101100100010000011;  // -882278991 1957873795
      9'h46: T=64'b1100101010110010011011111010101001110100010111111001110111010000;  // -894275670 1952423376
      9'h47: T=64'b1100100111111011111001010010011101110100000010110101001111111010;  // -906238681 1946899450
      9'h48: T=64'b1100100101000101110111111110110101110011101101011110101111010000;  // -918167571 1941302224
      9'h49: T=64'b1100100010010000011000011011101001110011010111110110011000100101;  // -930061894 1935631909
      9'h4a: T=64'b1100011111011011011011000101000001110011000001111100001111001111;  // -941921200 1929888719
      9'h4b: T=64'b1100011100100111000000010110110101110010101011110000010110100110;  // -953745043 1924072870
      9'h4c: T=64'b1100011001110011001000101100111001110010010101010010110010000100;  // -965532978 1918184580
      9'h4d: T=64'b1100010110111111110100100010111101110001111110100011100101001000;  // -977284561 1912224072
      9'h4e: T=64'b1100010100001101000100010100100101110001100111100010110011010001;  // -988999351 1906191569
      9'h4f: T=64'b1100010001011010111000011101011101110001010000010000100000000100;  // -1000676905 1900087300
      9'h50: T=64'b1100001110101001010001011001000001110000111000101100101111000101;  // -1012316784 1893911493
      9'h51: T=64'b1100001011111000001111100010101101110000100000110111100011111110;  // -1023918549 1887664382
      9'h52: T=64'b1100001001000111110011010101101101110000001000110001000010011001;  // -1035481765 1881346201
      9'h53: T=64'b1100000110010111111101001101010001101111110000011001001110000100;  // -1047005996 1874957188
      9'h54: T=64'b1100000011101000101101100100100101101111010111110000001010110001;  // -1058490807 1868497585
      9'h55: T=64'b1100000000111010000100110110100101101110111110110101111100010001;  // -1069935767 1861967633
      9'h56: T=64'b1011111110001100000011011110001101101110100101101010100110011100;  // -1081340445 1855367580
      9'h57: T=64'b1011111011011110101001110110011001101110001100001110001101001001;  // -1092704410 1848697673
      9'h58: T=64'b1011111000110001111000011001110001101101110010100000110100010100;  // -1104027236 1841958164
      9'h59: T=64'b1011110110000101101111100011000001101101011000100010011111111001;  // -1115308496 1835149305
      9'h5a: T=64'b1011110011011010001111101100101101101100111110010011010011111011;  // -1126547765 1828271355
      9'h5b: T=64'b1011110000101111011001010001010001101100100011110011010100011011;  // -1137744620 1821324571
      9'h5c: T=64'b1011101110000101001100101011000001101100001001000010100101011111;  // -1148898640 1814309215
      9'h5d: T=64'b1011101011011011101010010100010001101011101110000001001011010000;  // -1160009404 1807225552
      9'h5e: T=64'b1011101000110010110010100111000101101011010010101111001001111000;  // -1171076495 1800073848
      9'h5f: T=64'b1011100110001010100101111101100101101010110111001100100101100100;  // -1182099495 1792854372
      9'h60: T=64'b1011100011100011000100110001101001101010011011011001100010100011;  // -1193077990 1785567395
      9'h61: T=64'b1011100000111100001111011101001001101001111111010110000101001010;  // -1204011566 1778213194
      9'h62: T=64'b1011011110010110000110011001110001101001100011000010010001101011;  // -1214899812 1770792043
      9'h63: T=64'b1011011011110000101010000001001001101001000110011110001100011111;  // -1225742318 1763304223
      9'h64: T=64'b1011011001001011111010101100110101101000101001101001111010000000;  // -1236538675 1755750016
      9'h65: T=64'b1011010110100111111000110110001101101000001100100101011110101010;  // -1247288477 1748129706
      9'h66: T=64'b1011010100000100100100110110100101100111101111010000111110111100;  // -1257991319 1740443580
      9'h67: T=64'b1011010001100001111111000111000101100111010001101100011111010111;  // -1268646799 1732691927
      9'h68: T=64'b1011001111000000001000000000110101100110110011111000000100011111;  // -1279254515 1724875039
      9'h69: T=64'b1011001100011110111111111100110001100110010101110011110010111011;  // -1289814068 1716993211
      9'h6a: T=64'b1011001001111110100111010011110101100101110111011111101111010010;  // -1300325059 1709046738
      9'h6b: T=64'b1011000111011110111110011110100101100101011000111011111110010001;  // -1310787095 1701035921
      9'h6c: T=64'b1011000101000000000101110101110001100100111010001000100100100101;  // -1321199780 1692961061
      9'h6d: T=64'b1011000010100001111101110001111001100100011011000101100110111111;  // -1331562722 1684822463
      9'h6e: T=64'b1011000000000100100110101011010001100011111011110011001010001111;  // -1341875532 1676620431
      9'h6f: T=64'b1010111101101000000000111010001001100011011100010001010011001100;  // -1352137822 1668355276
      9'h70: T=64'b1010111011001100001100110110110001100010111100100000000110101100;  // -1362349204 1660027308
      9'h71: T=64'b1010111000110001001010111001001001100010011100011111101001101000;  // -1372509294 1651636840
      9'h72: T=64'b1010110110010110111011011001001001100001111100010000000000111110;  // -1382617710 1643184190
      9'h73: T=64'b1010110011111101011110101110100101100001011011110001010001101011;  // -1392674071 1634669675
      9'h74: T=64'b1010110001100100110101010001000101100000111011000011100000101111;  // -1402677999 1626093615
      9'h75: T=64'b1010101111001100111111011000001101100000011010000110110011001110;  // -1412629117 1617456334
      9'h76: T=64'b1010101100110101111101011011011001011111111000111011001110001101;  // -1422527050 1608758157
      9'h77: T=64'b1010101010011111101111110001111001011111010111100000110110110010;  // -1432371426 1599999410
      9'h78: T=64'b1010101000001010010110110010111001011110110101110111110010001001;  // -1442161874 1591180425
      9'h79: T=64'b1010100101110101110010110101011101011110010100000000000101011101;  // -1451898025 1582301533
      9'h7a: T=64'b1010100011100010000100010000011101011101110001111001110101111011;  // -1461579513 1573363067
      9'h7b: T=64'b1010100001001111001011011010101101011101001111100101001000110110;  // -1471205973 1564365366
      9'h7c: T=64'b1010011110111101001000101010110001011100101101000010000011011111;  // -1480777044 1555308767
      9'h7d: T=64'b1010011100101011111100010111010001011100001010010000101011001100;  // -1490292364 1546193612
      9'h7e: T=64'b1010011010011011100110110110100101011011100111010001000101010011;  // -1499751575 1537020243
      9'h7f: T=64'b1010011000001100001000011110111001011011000100000011010111001110;  // -1509154322 1527789006
      9'h80: T=64'b1010010101111101100001100110011101011010100000100111100110011001;  // -1518500249 1518500249
      9'h81: T=64'b1010010011101111110010100011001001011001111100111101111000010010;  // -1527789006 1509154322
      9'h82: T=64'b1010010001100010111011101010110101011001011001000110010010010111;  // -1537020243 1499751575
      9'h83: T=64'b1010001111010110111101010011010001011000110101000000111010001100;  // -1546193612 1490292364
      9'h84: T=64'b1010001101001011110111110010000101011000010000101101110101010100;  // -1555308767 1480777044
      9'h85: T=64'b1010001011000001101011011100101001010111101100001101001001010101;  // -1564365366 1471205973
      9'h86: T=64'b1010001000111000011000101000010101010111000111011110111011111001;  // -1573363067 1461579513
      9'h87: T=64'b1010000110101111111111101010001101010110100010100011010010101001;  // -1582301533 1451898025
      9'h88: T=64'b1010000100101000100000110111011101010101111101011010010011010010;  // -1591180425 1442161874
      9'h89: T=64'b1010000010100001111100100100111001010101011000000100000011100010;  // -1599999410 1432371426
      9'h8a: T=64'b1010000000011100010011000111001101010100110010100000101001001010;  // -1608758157 1422527050
      9'h8b: T=64'b1001111110010111100100110011001001010100001100110000001001111101;  // -1617456334 1412629117
      9'h8c: T=64'b1001111100010011110001111101000101010011100110110010101011101111;  // -1626093615 1402677999
      9'h8d: T=64'b1001111010010000111010111001010101010011000000101000010100010111;  // -1634669675 1392674071
      9'h8e: T=64'b1001111000001110111111111100001001010010011010010001001001101110;  // -1643184190 1382617710
      9'h8f: T=64'b1001110110001110000001011001100001010001110011101101010001101110;  // -1651636840 1372509294
      9'h90: T=64'b1001110100001101111111100101010001010001001100111100110010010100;  // -1660027308 1362349204
      9'h91: T=64'b1001110010001110111010110011010001010000100101111111110001011110;  // -1668355276 1352137822
      9'h92: T=64'b1001110000010000110011010111000101001111111110110110010101001100;  // -1676620431 1341875532
      9'h93: T=64'b1001101110010011101001100100000101001111010111100000100011100010;  // -1684822463 1331562722
      9'h94: T=64'b1001101100010111011101101101101101001110101111111110100010100100;  // -1692961061 1321199780
      9'h95: T=64'b1001101010011100010000000110111101001110001000010000011000010111;  // -1701035921 1310787095
      9'h96: T=64'b1001101000100010000001000010111001001101100000010110001011000011;  // -1709046738 1300325059
      9'h97: T=64'b1001100110101000110000110100010101001100111000010000000000110100;  // -1716993211 1289814068
      9'h98: T=64'b1001100100110000011111101110000101001100001111111101111111110011;  // -1724875039 1279254515
      9'h99: T=64'b1001100010111001001110000010100101001011100111100000001110001111;  // -1732691927 1268646799
      9'h9a: T=64'b1001100001000010111100000100010001001010111110110110110010010111;  // -1740443580 1257991319
      9'h9b: T=64'b1001011111001101101010000101011001001010010110000001110010011101;  // -1748129706 1247288477
      9'h9c: T=64'b1001011101011001011000011000000001001001101101000001010100110011;  // -1755750016 1236538675
      9'h9d: T=64'b1001011011100110000111001110000101001001000011110101011111101110;  // -1763304223 1225742318
      9'h9e: T=64'b1001011001110011110110111001010101001000011010011110011001100100;  // -1770792043 1214899812
      9'h9f: T=64'b1001011000000010100111101011011001000111110000111100001000101110;  // -1778213194 1204011566
      9'ha0: T=64'b1001010110010010011001110101110101000111000111001110110011100110;  // -1785567395 1193077990
      9'ha1: T=64'b1001010100100011001101101001110001000110011101010110100000100111;  // -1792854372 1182099495
      9'ha2: T=64'b1001010010110101000011011000100001000101110011010011010110001111;  // -1800073848 1171076495
      9'ha3: T=64'b1001010001000111111011010011000001000101001001000101011010111100;  // -1807225552 1160009404
      9'ha4: T=64'b1001001111011011110101101010000101000100011110101100110101010000;  // -1814309215 1148898640
      9'ha5: T=64'b1001001101110000110010101110010101000011110100001001101011101100;  // -1821324571 1137744620
      9'ha6: T=64'b1001001100000110110010110000010101000011001001011100000100110101;  // -1828271355 1126547765
      9'ha7: T=64'b1001001010011101110110000000011101000010011110100100000111010000;  // -1835149305 1115308496
      9'ha8: T=64'b1001001000110101111100101110110001000001110011100001111001100100;  // -1841958164 1104027236
      9'ha9: T=64'b1001000111001111000111001011011101000001001000010101100010011010;  // -1848697673 1092704410
      9'haa: T=64'b1001000101101001010101100110010001000000011100111111001000011101;  // -1855367580 1081340445
      9'hab: T=64'b1001000100000100101000001110111100111111110001011110110010010111;  // -1861967633 1069935767
      9'hac: T=64'b1001000010100000111111010100111100111111000101110100100110110111;  // -1868497585 1058490807
      9'had: T=64'b1001000000111110011011000111110000111110011010000000101100101100;  // -1874957188 1047005996
      9'hae: T=64'b1000111111011100111011110110011100111101101110000011001010100101;  // -1881346201 1035481765
      9'haf: T=64'b1000111101111100100001110000001000111101000001111100000111010101;  // -1887664382 1023918549
      9'hb0: T=64'b1000111100011101001101000011101100111100010101101011101001110000;  // -1893911493 1012316784
      9'hb1: T=64'b1000111010111110111101111111110000111011101001010001111000101001;  // -1900087300 1000676905
      9'hb2: T=64'b1000111001100001110100110010111100111010111100101110111010110111;  // -1906191569 988999351
      9'hb3: T=64'b1000111000000101110001101011100000111010010000000010110111010001;  // -1912224072 977284561
      9'hb4: T=64'b1000110110101010110100110111110000111001100011001101110100110010;  // -1918184580 965532978
      9'hb5: T=64'b1000110101010000111110100101101000111000110110001111111010010011;  // -1924072870 953745043
      9'hb6: T=64'b1000110011111000001111000011000100111000001001001001001110110000;  // -1929888719 941921200
      9'hb7: T=64'b1000110010100000100110011101101100110111011011111001111001000110;  // -1935631909 930061894
      9'hb8: T=64'b1000110001001010000101000011000000110110101110100010000000010011;  // -1941302224 918167571
      9'hb9: T=64'b1000101111110100101011000000011000110110000001000001101011011001;  // -1946899450 906238681
      9'hba: T=64'b1000101110100000011000100011000000110101010011011001000001010110;  // -1952423376 894275670
      9'hbb: T=64'b1000101101001101001101110111110100110100100101101000001001001111;  // -1957873795 882278991
      9'hbc: T=64'b1000101011111011001011001011110000110011110111101111001010000111;  // -1963250500 870249095
      9'hbd: T=64'b1000101010101010010000101011010100110011001001101110001011000010;  // -1968553291 858186434
      9'hbe: T=64'b1000101001011010011110100011001000110010011011100101010011000111;  // -1973781966 846091463
      9'hbf: T=64'b1000101000001011110100111111011000110001101101010100101001011101;  // -1978936330 833964637
      9'hc0: T=64'b1000100110111110010100001100010000110000111110111100010101001101;  // -1984016188 821806413
      9'hc1: T=64'b1000100101110001111100010101101100110000010000011100011101100000;  // -1989021349 809617248
      9'hc2: T=64'b1000100100100110101101100111100000101111100001110101001001100010;  // -1993951624 797397602
      9'hc3: T=64'b1000100011011100101000001101010000101110110011000110100000011110;  // -1998806828 785147934
      9'hc4: T=64'b1000100010010011101100010010011000101110000100010000101001100010;  // -2003586778 772868706
      9'hc5: T=64'b1000100001001011111010000010000100101101010101010011101011111011;  // -2008291295 760560379
      9'hc6: T=64'b1000100000000101010001100111100000101100100110001111101110111010;  // -2012920200 748223418
      9'hc7: T=64'b1000011110111111110011001101100000101011110111000100111001101111;  // -2017473320 735858287
      9'hc8: T=64'b1000011101111011011110111110110100101011000111110011010011101011;  // -2021950483 723465451
      9'hc9: T=64'b1000011100111000010101000101111100101010011000011011000100000001;  // -2026351521 711045377
      9'hca: T=64'b1000011011110110010101101101010000101001101000111100010010000101;  // -2030676268 698598533
      9'hcb: T=64'b1000011010110101100000111110111100101000111001010111000101001010;  // -2034924561 686125386
      9'hcc: T=64'b1000011001110101110111000101000000101000001001101011100100101000;  // -2039096240 673626408
      9'hcd: T=64'b1000011000110111011000001001001100100111011001111001110111110100;  // -2043191149 661102068
      9'hce: T=64'b1000010111111010000100010101010000100110101010000010000110000101;  // -2047209132 648552837
      9'hcf: T=64'b1000010110111101111011110010100000100101111010000100010110110110;  // -2051150040 635979190
      9'hd0: T=64'b1000010110000010111110101010011000100101001010000000110001011101;  // -2055013722 623381597
      9'hd1: T=64'b1000010101001001001101000101110100100100011001110111011101010111;  // -2058800035 610760535
      9'hd2: T=64'b1000010100010000100111001101110100100011101001101000100001111110;  // -2062508835 598116478
      9'hd3: T=64'b1000010011011001001101001011001000100010111001010100000110101111;  // -2066139982 585449903
      9'hd4: T=64'b1000010010100010111111000110001100100010001000111010010011000101;  // -2069693341 572761285
      9'hd5: T=64'b1000010001101101111101000111100000100001011000011011001110011111;  // -2073168776 560051103
      9'hd6: T=64'b1000010000111010000111010111000100100000100111110111000000011100;  // -2076566159 547319836
      9'hd7: T=64'b1000010000000111011101111101000100011111110111001101110000011011;  // -2079885359 534567963
      9'hd8: T=64'b1000001111010110000001000001001100011111000110011111100101111011;  // -2083126253 521795963
      9'hd9: T=64'b1000001110100101110000101011000100011110010101101100101000011110;  // -2086288719 509004318
      9'hda: T=64'b1000001101110110101101000010001100011101100100110100111111100101;  // -2089372637 496193509
      9'hdb: T=64'b1000001101001000110110001101110100011100110011111000110010110011;  // -2092377891 483364019
      9'hdc: T=64'b1000001100011100001100010100111100011100000010111000001001101010;  // -2095304369 470516330
      9'hdd: T=64'b1000001011110000101111011110100100011011010001110011001011101111;  // -2098151959 457650927
      9'hde: T=64'b1000001011000110011111110001010100011010100000101010000000100101;  // -2100920555 444768293
      9'hdf: T=64'b1000001010011101011101010011101100011001101111011100101111110011;  // -2103610053 431868915
      9'he0: T=64'b1000001001110101101000001100000100011000111110001011100000111100;  // -2106220351 418953276
      9'he1: T=64'b1000001001001111000000100000100100011000001100110110011011101000;  // -2108751351 406021864
      9'he2: T=64'b1000001000101001100110010111001000010111011011011101100111011110;  // -2111202958 393075166
      9'he3: T=64'b1000001000000101011001110101100100010110101010000001001100000101;  // -2113575079 380113669
      9'he4: T=64'b1000000111100010011011000001011100010101111000100001010001000100;  // -2115867625 367137860
      9'he5: T=64'b1000000111000000101010000000001000010101000110111101111110000101;  // -2118080510 354148229
      9'he6: T=64'b1000000110100000000110110110111000010100010101010111011010110001;  // -2120213650 341145265
      9'he7: T=64'b1000000110000000110001101010101000010011100011101101101110110001;  // -2122266966 328129457
      9'he8: T=64'b1000000101100010101010100000010100010010110010000001000001101110;  // -2124240379 315101294
      9'he9: T=64'b1000000101000101110001011100100000010010000000010001011011010101;  // -2126133816 302061269
      9'hea: T=64'b1000000100101010000110100011101100010001001110011111000011001111;  // -2127947205 289009871
      9'heb: T=64'b1000000100001111101001111010000100010000011100101010000001001000;  // -2129680479 275947592
      9'hec: T=64'b1000000011110110011011100011110100001111101010110010011100101011;  // -2131333571 262874923
      9'hed: T=64'b1000000011011110011011100100110100001110111000111000011101100110;  // -2132906419 249792358
      9'hee: T=64'b1000000011000111101010000000101100001110000110111100001011100100;  // -2134398965 236700388
      9'hef: T=64'b1000000010110010000110111011000000001101010100111101101110010010;  // -2135811152 223599506
      9'hf0: T=64'b1000000010011101110010010111001000001100100010111101001101011110;  // -2137142926 210490206
      9'hf1: T=64'b1000000010001010101100011000000100001011110000111010110000110101;  // -2138394239 197372981
      9'hf2: T=64'b1000000001111000110101000000111000001010111110110110100000000101;  // -2139565042 184248325
      9'hf3: T=64'b1000000001101000001100010100010000001010001100110000100010111100;  // -2140655292 171116732
      9'hf4: T=64'b1000000001011000110010010100110100001001011010101001000001001001;  // -2141664947 157978697
      9'hf5: T=64'b1000000001001010100111000100111000001000101000100000000010011010;  // -2142593970 144834714
      9'hf6: T=64'b1000000000111101101010100110101100000111110110010101101110011110;  // -2143442325 131685278
      9'hf7: T=64'b1000000000110001111100111100001100000111000100001010001101000101;  // -2144209981 118530885
      9'hf8: T=64'b1000000000100111011110000111001100000110010001111101100101111100;  // -2144896909 105372028
      9'hf9: T=64'b1000000000011110001110001001011000000101011111110000000000110101;  // -2145503082 92209205
      9'hfa: T=64'b1000000000010110001101000100000100000100101101100001100101011101;  // -2146028479 79042909
      9'hfb: T=64'b1000000000001111011010111000100100000011111011010010011011100110;  // -2146473079 65873638
      9'hfc: T=64'b1000000000001001110111100111111100000011001001000010101010111111;  // -2146836865 52701887
      9'hfd: T=64'b1000000000000101100011010011000000000010010110110010011011010111;  // -2147119824 39528151
      9'hfe: T=64'b1000000000000010011101111010011100000001100100100001110100100000;  // -2147321945 26352928
      9'hff: T=64'b1000000000000000100111011110101100000000110010010000111110001000;  // -2147443221 13176712
      9'h100: T=64'b1000000000000000000000000000000100000000000000000000000000000000;  // -2147483647     0
      9'h101: T=64'b1000000000000000100111011110101111111111001101101111000001111000;  // -2147443221 -13176712
      9'h102: T=64'b1000000000000010011101111010011111111110011011011110001011100000;  // -2147321945 -26352928
      9'h103: T=64'b1000000000000101100011010011000011111101101001001101100100101001;  // -2147119824 -39528151
      9'h104: T=64'b1000000000001001110111100111111111111100110110111101010101000001;  // -2146836865 -52701887
      9'h105: T=64'b1000000000001111011010111000100111111100000100101101100100011010;  // -2146473079 -65873638
      9'h106: T=64'b1000000000010110001101000100000111111011010010011110011010100011;  // -2146028479 -79042909
      9'h107: T=64'b1000000000011110001110001001011011111010100000001111111111001011;  // -2145503082 -92209205
      9'h108: T=64'b1000000000100111011110000111001111111001101110000010011010000100;  // -2144896909 -105372028
      9'h109: T=64'b1000000000110001111100111100001111111000111011110101110010111011;  // -2144209981 -118530885
      9'h10a: T=64'b1000000000111101101010100110101111111000001001101010010001100010;  // -2143442325 -131685278
      9'h10b: T=64'b1000000001001010100111000100111011110111010111011111111101100110;  // -2142593970 -144834714
      9'h10c: T=64'b1000000001011000110010010100110111110110100101010110111110110111;  // -2141664947 -157978697
      9'h10d: T=64'b1000000001101000001100010100010011110101110011001111011101000100;  // -2140655292 -171116732
      9'h10e: T=64'b1000000001111000110101000000111011110101000001001001011111111011;  // -2139565042 -184248325
      9'h10f: T=64'b1000000010001010101100011000000111110100001111000101001111001011;  // -2138394239 -197372981
      9'h110: T=64'b1000000010011101110010010111001011110011011101000010110010100010;  // -2137142926 -210490206
      9'h111: T=64'b1000000010110010000110111011000011110010101011000010010001101110;  // -2135811152 -223599506
      9'h112: T=64'b1000000011000111101010000000101111110001111001000011110100011100;  // -2134398965 -236700388
      9'h113: T=64'b1000000011011110011011100100110111110001000111000111100010011010;  // -2132906419 -249792358
      9'h114: T=64'b1000000011110110011011100011110111110000010101001101100011010101;  // -2131333571 -262874923
      9'h115: T=64'b1000000100001111101001111010000111101111100011010101111110111000;  // -2129680479 -275947592
      9'h116: T=64'b1000000100101010000110100011101111101110110001100000111100110001;  // -2127947205 -289009871
      9'h117: T=64'b1000000101000101110001011100100011101101111111101110100100101011;  // -2126133816 -302061269
      9'h118: T=64'b1000000101100010101010100000010111101101001101111110111110010010;  // -2124240379 -315101294
      9'h119: T=64'b1000000110000000110001101010101011101100011100010010010001001111;  // -2122266966 -328129457
      9'h11a: T=64'b1000000110100000000110110110111011101011101010101000100101001111;  // -2120213650 -341145265
      9'h11b: T=64'b1000000111000000101010000000001011101010111001000010000001111011;  // -2118080510 -354148229
      9'h11c: T=64'b1000000111100010011011000001011111101010000111011110101110111100;  // -2115867625 -367137860
      9'h11d: T=64'b1000001000000101011001110101100111101001010101111110110011111011;  // -2113575079 -380113669
      9'h11e: T=64'b1000001000101001100110010111001011101000100100100010011000100010;  // -2111202958 -393075166
      9'h11f: T=64'b1000001001001111000000100000100111100111110011001001100100011000;  // -2108751351 -406021864
      9'h120: T=64'b1000001001110101101000001100000111100111000001110100011111000100;  // -2106220351 -418953276
      9'h121: T=64'b1000001010011101011101010011101111100110010000100011010000001101;  // -2103610053 -431868915
      9'h122: T=64'b1000001011000110011111110001010111100101011111010101111111011011;  // -2100920555 -444768293
      9'h123: T=64'b1000001011110000101111011110100111100100101110001100110100010001;  // -2098151959 -457650927
      9'h124: T=64'b1000001100011100001100010100111111100011111101000111110110010110;  // -2095304369 -470516330
      9'h125: T=64'b1000001101001000110110001101110111100011001100000111001101001101;  // -2092377891 -483364019
      9'h126: T=64'b1000001101110110101101000010001111100010011011001011000000011011;  // -2089372637 -496193509
      9'h127: T=64'b1000001110100101110000101011000111100001101010010011010111100010;  // -2086288719 -509004318
      9'h128: T=64'b1000001111010110000001000001001111100000111001100000011010000101;  // -2083126253 -521795963
      9'h129: T=64'b1000010000000111011101111101000111100000001000110010001111100101;  // -2079885359 -534567963
      9'h12a: T=64'b1000010000111010000111010111000111011111011000001000111111100100;  // -2076566159 -547319836
      9'h12b: T=64'b1000010001101101111101000111100011011110100111100100110001100001;  // -2073168776 -560051103
      9'h12c: T=64'b1000010010100010111111000110001111011101110111000101101100111011;  // -2069693341 -572761285
      9'h12d: T=64'b1000010011011001001101001011001011011101000110101011111001010001;  // -2066139982 -585449903
      9'h12e: T=64'b1000010100010000100111001101110111011100010110010111011110000010;  // -2062508835 -598116478
      9'h12f: T=64'b1000010101001001001101000101110111011011100110001000100010101001;  // -2058800035 -610760535
      9'h130: T=64'b1000010110000010111110101010011011011010110101111111001110100011;  // -2055013722 -623381597
      9'h131: T=64'b1000010110111101111011110010100011011010000101111011101001001010;  // -2051150040 -635979190
      9'h132: T=64'b1000010111111010000100010101010011011001010101111101111001111011;  // -2047209132 -648552837
      9'h133: T=64'b1000011000110111011000001001001111011000100110000110001000001100;  // -2043191149 -661102068
      9'h134: T=64'b1000011001110101110111000101000011010111110110010100011011011000;  // -2039096240 -673626408
      9'h135: T=64'b1000011010110101100000111110111111010111000110101000111010110110;  // -2034924561 -686125386
      9'h136: T=64'b1000011011110110010101101101010011010110010111000011101101111011;  // -2030676268 -698598533
      9'h137: T=64'b1000011100111000010101000101111111010101100111100100111011111111;  // -2026351521 -711045377
      9'h138: T=64'b1000011101111011011110111110110111010100111000001100101100010101;  // -2021950483 -723465451
      9'h139: T=64'b1000011110111111110011001101100011010100001000111011000110010001;  // -2017473320 -735858287
      9'h13a: T=64'b1000100000000101010001100111100011010011011001110000010001000110;  // -2012920200 -748223418
      9'h13b: T=64'b1000100001001011111010000010000111010010101010101100010100000101;  // -2008291295 -760560379
      9'h13c: T=64'b1000100010010011101100010010011011010001111011101111010110011110;  // -2003586778 -772868706
      9'h13d: T=64'b1000100011011100101000001101010011010001001100111001011111100010;  // -1998806828 -785147934
      9'h13e: T=64'b1000100100100110101101100111100011010000011110001010110110011110;  // -1993951624 -797397602
      9'h13f: T=64'b1000100101110001111100010101101111001111101111100011100010100000;  // -1989021349 -809617248
      9'h140: T=64'b1000100110111110010100001100010011001111000001000011101010110011;  // -1984016188 -821806413
      9'h141: T=64'b1000101000001011110100111111011011001110010010101011010110100011;  // -1978936330 -833964637
      9'h142: T=64'b1000101001011010011110100011001011001101100100011010101100111001;  // -1973781966 -846091463
      9'h143: T=64'b1000101010101010010000101011010111001100110110010001110100111110;  // -1968553291 -858186434
      9'h144: T=64'b1000101011111011001011001011110011001100001000010000110101111001;  // -1963250500 -870249095
      9'h145: T=64'b1000101101001101001101110111110111001011011010010111110110110001;  // -1957873795 -882278991
      9'h146: T=64'b1000101110100000011000100011000011001010101100100110111110101010;  // -1952423376 -894275670
      9'h147: T=64'b1000101111110100101011000000011011001001111110111110010100100111;  // -1946899450 -906238681
      9'h148: T=64'b1000110001001010000101000011000011001001010001011101111111101101;  // -1941302224 -918167571
      9'h149: T=64'b1000110010100000100110011101101111001000100100000110000110111010;  // -1935631909 -930061894
      9'h14a: T=64'b1000110011111000001111000011000111000111110110110110110001010000;  // -1929888719 -941921200
      9'h14b: T=64'b1000110101010000111110100101101011000111001001110000000101101101;  // -1924072870 -953745043
      9'h14c: T=64'b1000110110101010110100110111110011000110011100110010001011001110;  // -1918184580 -965532978
      9'h14d: T=64'b1000111000000101110001101011100011000101101111111101001000101111;  // -1912224072 -977284561
      9'h14e: T=64'b1000111001100001110100110010111111000101000011010001000101001001;  // -1906191569 -988999351
      9'h14f: T=64'b1000111010111110111101111111110011000100010110101110000111010111;  // -1900087300 -1000676905
      9'h150: T=64'b1000111100011101001101000011101111000011101010010100010110010000;  // -1893911493 -1012316784
      9'h151: T=64'b1000111101111100100001110000001011000010111110000011111000101011;  // -1887664382 -1023918549
      9'h152: T=64'b1000111111011100111011110110011111000010010001111100110101011011;  // -1881346201 -1035481765
      9'h153: T=64'b1001000000111110011011000111110011000001100101111111010011010100;  // -1874957188 -1047005996
      9'h154: T=64'b1001000010100000111111010100111111000000111010001011011001001001;  // -1868497585 -1058490807
      9'h155: T=64'b1001000100000100101000001110111111000000001110100001001101101001;  // -1861967633 -1069935767
      9'h156: T=64'b1001000101101001010101100110010010111111100011000000110111100011;  // -1855367580 -1081340445
      9'h157: T=64'b1001000111001111000111001011011110111110110111101010011101100110;  // -1848697673 -1092704410
      9'h158: T=64'b1001001000110101111100101110110010111110001100011110000110011100;  // -1841958164 -1104027236
      9'h159: T=64'b1001001010011101110110000000011110111101100001011011111000110000;  // -1835149305 -1115308496
      9'h15a: T=64'b1001001100000110110010110000010110111100110110100011111011001011;  // -1828271355 -1126547765
      9'h15b: T=64'b1001001101110000110010101110010110111100001011110110010100010100;  // -1821324571 -1137744620
      9'h15c: T=64'b1001001111011011110101101010000110111011100001010011001010110000;  // -1814309215 -1148898640
      9'h15d: T=64'b1001010001000111111011010011000010111010110110111010100101000100;  // -1807225552 -1160009404
      9'h15e: T=64'b1001010010110101000011011000100010111010001100101100101001110001;  // -1800073848 -1171076495
      9'h15f: T=64'b1001010100100011001101101001110010111001100010101001011111011001;  // -1792854372 -1182099495
      9'h160: T=64'b1001010110010010011001110101110110111000111000110001001100011010;  // -1785567395 -1193077990
      9'h161: T=64'b1001011000000010100111101011011010111000001111000011110111010010;  // -1778213194 -1204011566
      9'h162: T=64'b1001011001110011110110111001010110110111100101100001100110011100;  // -1770792043 -1214899812
      9'h163: T=64'b1001011011100110000111001110000110110110111100001010100000010010;  // -1763304223 -1225742318
      9'h164: T=64'b1001011101011001011000011000000010110110010010111110101011001101;  // -1755750016 -1236538675
      9'h165: T=64'b1001011111001101101010000101011010110101101001111110001101100011;  // -1748129706 -1247288477
      9'h166: T=64'b1001100001000010111100000100010010110101000001001001001101101001;  // -1740443580 -1257991319
      9'h167: T=64'b1001100010111001001110000010100110110100011000011111110001110001;  // -1732691927 -1268646799
      9'h168: T=64'b1001100100110000011111101110000110110011110000000010000000001101;  // -1724875039 -1279254515
      9'h169: T=64'b1001100110101000110000110100010110110011000111101111111111001100;  // -1716993211 -1289814068
      9'h16a: T=64'b1001101000100010000001000010111010110010011111101001110100111101;  // -1709046738 -1300325059
      9'h16b: T=64'b1001101010011100010000000110111110110001110111101111100111101001;  // -1701035921 -1310787095
      9'h16c: T=64'b1001101100010111011101101101101110110001010000000001011101011100;  // -1692961061 -1321199780
      9'h16d: T=64'b1001101110010011101001100100000110110000101000011111011100011110;  // -1684822463 -1331562722
      9'h16e: T=64'b1001110000010000110011010111000110110000000001001001101010110100;  // -1676620431 -1341875532
      9'h16f: T=64'b1001110010001110111010110011010010101111011010000000001110100010;  // -1668355276 -1352137822
      9'h170: T=64'b1001110100001101111111100101010010101110110011000011001101101100;  // -1660027308 -1362349204
      9'h171: T=64'b1001110110001110000001011001100010101110001100010010101110010010;  // -1651636840 -1372509294
      9'h172: T=64'b1001111000001110111111111100001010101101100101101110110110010010;  // -1643184190 -1382617710
      9'h173: T=64'b1001111010010000111010111001010110101100111111010111101011101001;  // -1634669675 -1392674071
      9'h174: T=64'b1001111100010011110001111101000110101100011001001101010100010001;  // -1626093615 -1402677999
      9'h175: T=64'b1001111110010111100100110011001010101011110011001111110110000011;  // -1617456334 -1412629117
      9'h176: T=64'b1010000000011100010011000111001110101011001101011111010110110110;  // -1608758157 -1422527050
      9'h177: T=64'b1010000010100001111100100100111010101010100111111011111100011110;  // -1599999410 -1432371426
      9'h178: T=64'b1010000100101000100000110111011110101010000010100101101100101110;  // -1591180425 -1442161874
      9'h179: T=64'b1010000110101111111111101010001110101001011101011100101101010111;  // -1582301533 -1451898025
      9'h17a: T=64'b1010001000111000011000101000010110101000111000100001000100000111;  // -1573363067 -1461579513
      9'h17b: T=64'b1010001011000001101011011100101010101000010011110010110110101011;  // -1564365366 -1471205973
      9'h17c: T=64'b1010001101001011110111110010000110100111101111010010001010101100;  // -1555308767 -1480777044
      9'h17d: T=64'b1010001111010110111101010011010010100111001010111111000101110100;  // -1546193612 -1490292364
      9'h17e: T=64'b1010010001100010111011101010110110100110100110111001101101101001;  // -1537020243 -1499751575
      9'h17f: T=64'b1010010011101111110010100011001010100110000011000010000111101110;  // -1527789006 -1509154322
      9'h180: T=64'b1010010101111101100001100110011110100101011111011000011001100111;  // -1518500249 -1518500249
      9'h181: T=64'b1010011000001100001000011110111010100100111011111100101000110010;  // -1509154322 -1527789006
      9'h182: T=64'b1010011010011011100110110110100110100100011000101110111010101101;  // -1499751575 -1537020243
      9'h183: T=64'b1010011100101011111100010111010010100011110101101111010100110100;  // -1490292364 -1546193612
      9'h184: T=64'b1010011110111101001000101010110010100011010010111101111100100001;  // -1480777044 -1555308767
      9'h185: T=64'b1010100001001111001011011010101110100010110000011010110111001010;  // -1471205973 -1564365366
      9'h186: T=64'b1010100011100010000100010000011110100010001110000110001010000101;  // -1461579513 -1573363067
      9'h187: T=64'b1010100101110101110010110101011110100001101011111111111010100011;  // -1451898025 -1582301533
      9'h188: T=64'b1010101000001010010110110010111010100001001010001000001101110111;  // -1442161874 -1591180425
      9'h189: T=64'b1010101010011111101111110001111010100000101000011111001001001110;  // -1432371426 -1599999410
      9'h18a: T=64'b1010101100110101111101011011011010100000000111000100110001110011;  // -1422527050 -1608758157
      9'h18b: T=64'b1010101111001100111111011000001110011111100101111001001100110010;  // -1412629117 -1617456334
      9'h18c: T=64'b1010110001100100110101010001000110011111000100111100011111010001;  // -1402677999 -1626093615
      9'h18d: T=64'b1010110011111101011110101110100110011110100100001110101110010101;  // -1392674071 -1634669675
      9'h18e: T=64'b1010110110010110111011011001001010011110000011101111111111000010;  // -1382617710 -1643184190
      9'h18f: T=64'b1010111000110001001010111001001010011101100011100000010110011000;  // -1372509294 -1651636840
      9'h190: T=64'b1010111011001100001100110110110010011101000011011111111001010100;  // -1362349204 -1660027308
      9'h191: T=64'b1010111101101000000000111010001010011100100011101110101100110100;  // -1352137822 -1668355276
      9'h192: T=64'b1011000000000100100110101011010010011100000100001100110101110001;  // -1341875532 -1676620431
      9'h193: T=64'b1011000010100001111101110001111010011011100100111010011001000001;  // -1331562722 -1684822463
      9'h194: T=64'b1011000101000000000101110101110010011011000101110111011011011011;  // -1321199780 -1692961061
      9'h195: T=64'b1011000111011110111110011110100110011010100111000100000001101111;  // -1310787095 -1701035921
      9'h196: T=64'b1011001001111110100111010011110110011010001000100000010000101110;  // -1300325059 -1709046738
      9'h197: T=64'b1011001100011110111111111100110010011001101010001100001101000101;  // -1289814068 -1716993211
      9'h198: T=64'b1011001111000000001000000000110110011001001100000111111011100001;  // -1279254515 -1724875039
      9'h199: T=64'b1011010001100001111111000111000110011000101110010011100000101001;  // -1268646799 -1732691927
      9'h19a: T=64'b1011010100000100100100110110100110011000010000101111000001000100;  // -1257991319 -1740443580
      9'h19b: T=64'b1011010110100111111000110110001110010111110011011010100001010110;  // -1247288477 -1748129706
      9'h19c: T=64'b1011011001001011111010101100110110010111010110010110000110000000;  // -1236538675 -1755750016
      9'h19d: T=64'b1011011011110000101010000001001010010110111001100001110011100001;  // -1225742318 -1763304223
      9'h19e: T=64'b1011011110010110000110011001110010010110011100111101101110010101;  // -1214899812 -1770792043
      9'h19f: T=64'b1011100000111100001111011101001010010110000000101001111010110110;  // -1204011566 -1778213194
      9'h1a0: T=64'b1011100011100011000100110001101010010101100100100110011101011101;  // -1193077990 -1785567395
      9'h1a1: T=64'b1011100110001010100101111101100110010101001000110011011010011100;  // -1182099495 -1792854372
      9'h1a2: T=64'b1011101000110010110010100111000110010100101101010000110110001000;  // -1171076495 -1800073848
      9'h1a3: T=64'b1011101011011011101010010100010010010100010001111110110100110000;  // -1160009404 -1807225552
      9'h1a4: T=64'b1011101110000101001100101011000010010011110110111101011010100001;  // -1148898640 -1814309215
      9'h1a5: T=64'b1011110000101111011001010001010010010011011100001100101011100101;  // -1137744620 -1821324571
      9'h1a6: T=64'b1011110011011010001111101100101110010011000001101100101100000101;  // -1126547765 -1828271355
      9'h1a7: T=64'b1011110110000101101111100011000010010010100111011101100000000111;  // -1115308496 -1835149305
      9'h1a8: T=64'b1011111000110001111000011001110010010010001101011111001011101100;  // -1104027236 -1841958164
      9'h1a9: T=64'b1011111011011110101001110110011010010001110011110001110010110111;  // -1092704410 -1848697673
      9'h1aa: T=64'b1011111110001100000011011110001110010001011010010101011001100100;  // -1081340445 -1855367580
      9'h1ab: T=64'b1100000000111010000100110110100110010001000001001010000011101111;  // -1069935767 -1861967633
      9'h1ac: T=64'b1100000011101000101101100100100110010000101000001111110101001111;  // -1058490807 -1868497585
      9'h1ad: T=64'b1100000110010111111101001101010010010000001111100110110001111100;  // -1047005996 -1874957188
      9'h1ae: T=64'b1100001001000111110011010101101110001111110111001110111101100111;  // -1035481765 -1881346201
      9'h1af: T=64'b1100001011111000001111100010101110001111011111001000011100000010;  // -1023918549 -1887664382
      9'h1b0: T=64'b1100001110101001010001011001000010001111000111010011010000111011;  // -1012316784 -1893911493
      9'h1b1: T=64'b1100010001011010111000011101011110001110101111101111011111111100;  // -1000676905 -1900087300
      9'h1b2: T=64'b1100010100001101000100010100100110001110011000011101001100101111;  // -988999351 -1906191569
      9'h1b3: T=64'b1100010110111111110100100010111110001110000001011100011010111000;  // -977284561 -1912224072
      9'h1b4: T=64'b1100011001110011001000101100111010001101101010101101001101111100;  // -965532978 -1918184580
      9'h1b5: T=64'b1100011100100111000000010110110110001101010100001111101001011010;  // -953745043 -1924072870
      9'h1b6: T=64'b1100011111011011011011000101000010001100111110000011110000110001;  // -941921200 -1929888719
      9'h1b7: T=64'b1100100010010000011000011011101010001100101000001001100111011011;  // -930061894 -1935631909
      9'h1b8: T=64'b1100100101000101110111111110110110001100010010100001010000110000;  // -918167571 -1941302224
      9'h1b9: T=64'b1100100111111011111001010010011110001011111101001010110000000110;  // -906238681 -1946899450
      9'h1ba: T=64'b1100101010110010011011111010101010001011101000000110001000110000;  // -894275670 -1952423376
      9'h1bb: T=64'b1100101101101001011111011011000110001011010011010011011101111101;  // -882278991 -1957873795
      9'h1bc: T=64'b1100110000100001000011010111100110001010111110110010110010111100;  // -870249095 -1963250500
      9'h1bd: T=64'b1100110011011001000111010011111010001010101010100100001010110101;  // -858186434 -1968553291
      9'h1be: T=64'b1100110110010001101010110011100110001010010110100111101000110010;  // -846091463 -1973781966
      9'h1bf: T=64'b1100111001001010101101011010001110001010000010111101001111110110;  // -833964637 -1978936330
      9'h1c0: T=64'b1100111100000100001110101011001110001001101111100101000011000100;  // -821806413 -1984016188
      9'h1c1: T=64'b1100111110111110001110001010000010001001011100011111000101011011;  // -809617248 -1989021349
      9'h1c2: T=64'b1101000001111000101011011001111010001001001001101011011001111000;  // -797397602 -1993951624
      9'h1c3: T=64'b1101000100110011100101111110001010001000110111001010000011010100;  // -785147934 -1998806828
      9'h1c4: T=64'b1101000111101110111101011001111010001000100100111011000100100110;  // -772868706 -2003586778
      9'h1c5: T=64'b1101001010101010110001010000010110001000010010111110100000100001;  // -760560379 -2008291295
      9'h1c6: T=64'b1101001101100111000001000100011010001000000001010100011001111000;  // -748223418 -2012920200
      9'h1c7: T=64'b1101010000100011101100011001000110000111101111111100110011011000;  // -735858287 -2017473320
      9'h1c8: T=64'b1101010011100000110010110001010110000111011110110111101111101101;  // -723465451 -2021950483
      9'h1c9: T=64'b1101010110011110010011101111111110000111001110000101010001011111;  // -711045377 -2026351521
      9'h1ca: T=64'b1101011001011100001110110111101110000110111101100101011011010100;  // -698598533 -2030676268
      9'h1cb: T=64'b1101011100011010100011101011011010000110101101011000001111101111;  // -686125386 -2034924561
      9'h1cc: T=64'b1101011111011001010001101101100010000110011101011101110001010000;  // -673626408 -2039096240
      9'h1cd: T=64'b1101100010011000011000100000110010000110001101110110000010010011;  // -661102068 -2043191149
      9'h1ce: T=64'b1101100101010111110111100111101110000101111110100001000101010100;  // -648552837 -2047209132
      9'h1cf: T=64'b1101101000010111101110100100101010000101101111011110111100101000;  // -635979190 -2051150040
      9'h1d0: T=64'b1101101011010111111100111010001110000101100000101111101010100110;  // -623381597 -2055013722
      9'h1d1: T=64'b1101101110011000100010001010100110000101010010010011010001011101;  // -610760535 -2058800035
      9'h1d2: T=64'b1101110001011001011101111000001010000101000100001001110011011101;  // -598116478 -2062508835
      9'h1d3: T=64'b1101110100011010101111100101000110000100110110010011010010110010;  // -585449903 -2066139982
      9'h1d4: T=64'b1101110111011100010110110011101110000100101000101111110001100011;  // -572761285 -2069693341
      9'h1d5: T=64'b1101111010011110010011000110000110000100011011011111010001111000;  // -560051103 -2073168776
      9'h1d6: T=64'b1101111101100000100011111110010010000100001110100001110101110001;  // -547319836 -2076566159
      9'h1d7: T=64'b1110000000100011001000111110010110000100000001110111011111010001;  // -534567963 -2079885359
      9'h1d8: T=64'b1110000011100110000001101000010110000011110101100000010000010011;  // -521795963 -2083126253
      9'h1d9: T=64'b1110000110101001001101011110001010000011101001011100001010110001;  // -509004318 -2086288719
      9'h1da: T=64'b1110001001101100101100000001101110000011011101101011010000100011;  // -496193509 -2089372637
      9'h1db: T=64'b1110001100110000011100110100110110000011010010001101100011011101;  // -483364019 -2092377891
      9'h1dc: T=64'b1110001111110100011111011001011010000011000111000011000101001111;  // -470516330 -2095304369
      9'h1dd: T=64'b1110010010111000110011010001000110000010111100001011110111101001;  // -457650927 -2098151959
      9'h1de: T=64'b1110010101111101010111111101101110000010110001100111111100010101;  // -444768293 -2100920555
      9'h1df: T=64'b1110011001000010001101000000110110000010100111010111010100111011;  // -431868915 -2103610053
      9'h1e0: T=64'b1110011100000111010001111100010010000010011101011010000011000001;  // -418953276 -2106220351
      9'h1e1: T=64'b1110011111001100100110010001100010000010010011110000001000001001;  // -406021864 -2108751351
      9'h1e2: T=64'b1110100010010010001001100010001010000010001010011001100101110010;  // -393075166 -2111202958
      9'h1e3: T=64'b1110100101010111111011001111101110000010000001010110011101011001;  // -380113669 -2113575079
      9'h1e4: T=64'b1110101000011101111010111011110010000001111000100110110000010111;  // -367137860 -2115867625
      9'h1e5: T=64'b1110101011100100001000000111101110000001110000001010100000000010;  // -354148229 -2118080510
      9'h1e6: T=64'b1110101110101010100010010100111110000001101000000001101101101110;  // -341145265 -2120213650
      9'h1e7: T=64'b1110110001110001001001000100111110000001100000001100011010101010;  // -328129457 -2122266966
      9'h1e8: T=64'b1110110100110111111011111001001010000001011000101010101000000101;  // -315101294 -2124240379
      9'h1e9: T=64'b1110110111111110111010010010101110000001010001011100010111001000;  // -302061269 -2126133816
      9'h1ea: T=64'b1110111011000110000011110011000110000001001010100001101000111011;  // -289009871 -2127947205
      9'h1eb: T=64'b1110111110001101010111111011100010000001000011111010011110100001;  // -275947592 -2129680479
      9'h1ec: T=64'b1111000001010100110110001101010110000000111101100110111000111101;  // -262874923 -2131333571
      9'h1ed: T=64'b1111000100011100011110001001101010000000110111100110111001001101;  // -249792358 -2132906419
      9'h1ee: T=64'b1111000111100100001111010001110010000000110001111010100000001011;  // -236700388 -2134398965
      9'h1ef: T=64'b1111001010101100001001000110111010000000101100100001101110110000;  // -223599506 -2135811152
      9'h1f0: T=64'b1111001101110100001011001010001010000000100111011100100101110010;  // -210490206 -2137142926
      9'h1f1: T=64'b1111010000111100010100111100101110000000100010101011000110000001;  // -197372981 -2138394239
      9'h1f2: T=64'b1111010100000100100101111111101110000000011110001101010000001110;  // -184248325 -2139565042
      9'h1f3: T=64'b1111010111001100111101110100010010000000011010000011000101000100;  // -171116732 -2140655292
      9'h1f4: T=64'b1111011010010101011011111011011110000000010110001100100101001101;  // -157978697 -2141664947
      9'h1f5: T=64'b1111011101011101111111110110011010000000010010101001110001001110;  // -144834714 -2142593970
      9'h1f6: T=64'b1111100000100110101001000110001010000000001111011010101001101011;  // -131685278 -2143442325
      9'h1f7: T=64'b1111100011101111010111001011101110000000001100011111001111000011;  // -118530885 -2144209981
      9'h1f8: T=64'b1111100110111000001001101000010010000000001001110111100001110011;  // -105372028 -2144896909
      9'h1f9: T=64'b1111101010000000111111111100101110000000000111100011100010010110;  // -92209205 -2145503082
      9'h1fa: T=64'b1111101101001001111001101010001110000000000101100011010001000001;  // -79042909 -2146028479
      9'h1fb: T=64'b1111110000010010110110010001101010000000000011110110101110001001;  // -65873638 -2146473079
      9'h1fc: T=64'b1111110011011011110101010100000110000000000010011101111001111111;  // -52701887 -2146836865
      9'h1fd: T=64'b1111110110100100110110010010100110000000000001011000110100110000;  // -39528151 -2147119824
      9'h1fe: T=64'b1111111001101101111000101110000010000000000000100111011110100111;  // -26352928 -2147321945
      9'h1ff: T=64'b1111111100110110111100000111100010000000000000001001110111101011;  // -13176712 -2147443221
      default: T=64'b0;
    endcase

endmodule
