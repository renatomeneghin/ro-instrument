`timescale 1ns/10ps

module COREDDS_C0_COREDDS_C0_0_dds_qrtr_sin (index, sine);
  input  [8:0] index;
  output [17:0] sine;
  reg signed [17:0] sine/* synthesis syn_maxfan = 1000 */;

  always @ (index) 
    case (index) 
         0: sine = 18'b000000000000110010;  //         50 
         1: sine = 18'b000000000010010111;  //        151 
         2: sine = 18'b000000000011111011;  //        251 
         3: sine = 18'b000000000101100000;  //        352 
         4: sine = 18'b000000000111000100;  //        452 
         5: sine = 18'b000000001000101001;  //        553 
         6: sine = 18'b000000001010001101;  //        653 
         7: sine = 18'b000000001011110010;  //        754 
         8: sine = 18'b000000001101010110;  //        854 
         9: sine = 18'b000000001110111011;  //        955 
        10: sine = 18'b000000010000100000;  //       1056 
        11: sine = 18'b000000010010000100;  //       1156 
        12: sine = 18'b000000010011101001;  //       1257 
        13: sine = 18'b000000010101001101;  //       1357 
        14: sine = 18'b000000010110110010;  //       1458 
        15: sine = 18'b000000011000010110;  //       1558 
        16: sine = 18'b000000011001111011;  //       1659 
        17: sine = 18'b000000011011011111;  //       1759 
        18: sine = 18'b000000011101000100;  //       1860 
        19: sine = 18'b000000011110101000;  //       1960 
        20: sine = 18'b000000100000001101;  //       2061 
        21: sine = 18'b000000100001110001;  //       2161 
        22: sine = 18'b000000100011010101;  //       2261 
        23: sine = 18'b000000100100111010;  //       2362 
        24: sine = 18'b000000100110011110;  //       2462 
        25: sine = 18'b000000101000000011;  //       2563 
        26: sine = 18'b000000101001100111;  //       2663 
        27: sine = 18'b000000101011001100;  //       2764 
        28: sine = 18'b000000101100110000;  //       2864 
        29: sine = 18'b000000101110010101;  //       2965 
        30: sine = 18'b000000101111111001;  //       3065 
        31: sine = 18'b000000110001011101;  //       3165 
        32: sine = 18'b000000110011000010;  //       3266 
        33: sine = 18'b000000110100100110;  //       3366 
        34: sine = 18'b000000110110001011;  //       3467 
        35: sine = 18'b000000110111101111;  //       3567 
        36: sine = 18'b000000111001010011;  //       3667 
        37: sine = 18'b000000111010111000;  //       3768 
        38: sine = 18'b000000111100011100;  //       3868 
        39: sine = 18'b000000111110000001;  //       3969 
        40: sine = 18'b000000111111100101;  //       4069 
        41: sine = 18'b000001000001001001;  //       4169 
        42: sine = 18'b000001000010101110;  //       4270 
        43: sine = 18'b000001000100010010;  //       4370 
        44: sine = 18'b000001000101110110;  //       4470 
        45: sine = 18'b000001000111011010;  //       4570 
        46: sine = 18'b000001001000111111;  //       4671 
        47: sine = 18'b000001001010100011;  //       4771 
        48: sine = 18'b000001001100000111;  //       4871 
        49: sine = 18'b000001001101101100;  //       4972 
        50: sine = 18'b000001001111010000;  //       5072 
        51: sine = 18'b000001010000110100;  //       5172 
        52: sine = 18'b000001010010011000;  //       5272 
        53: sine = 18'b000001010011111100;  //       5372 
        54: sine = 18'b000001010101100001;  //       5473 
        55: sine = 18'b000001010111000101;  //       5573 
        56: sine = 18'b000001011000101001;  //       5673 
        57: sine = 18'b000001011010001101;  //       5773 
        58: sine = 18'b000001011011110001;  //       5873 
        59: sine = 18'b000001011101010101;  //       5973 
        60: sine = 18'b000001011110111001;  //       6073 
        61: sine = 18'b000001100000011101;  //       6173 
        62: sine = 18'b000001100010000010;  //       6274 
        63: sine = 18'b000001100011100110;  //       6374 
        64: sine = 18'b000001100101001010;  //       6474 
        65: sine = 18'b000001100110101110;  //       6574 
        66: sine = 18'b000001101000010010;  //       6674 
        67: sine = 18'b000001101001110110;  //       6774 
        68: sine = 18'b000001101011011010;  //       6874 
        69: sine = 18'b000001101100111110;  //       6974 
        70: sine = 18'b000001101110100010;  //       7074 
        71: sine = 18'b000001110000000110;  //       7174 
        72: sine = 18'b000001110001101001;  //       7273 
        73: sine = 18'b000001110011001101;  //       7373 
        74: sine = 18'b000001110100110001;  //       7473 
        75: sine = 18'b000001110110010101;  //       7573 
        76: sine = 18'b000001110111111001;  //       7673 
        77: sine = 18'b000001111001011101;  //       7773 
        78: sine = 18'b000001111011000001;  //       7873 
        79: sine = 18'b000001111100100100;  //       7972 
        80: sine = 18'b000001111110001000;  //       8072 
        81: sine = 18'b000001111111101100;  //       8172 
        82: sine = 18'b000010000001010000;  //       8272 
        83: sine = 18'b000010000010110011;  //       8371 
        84: sine = 18'b000010000100010111;  //       8471 
        85: sine = 18'b000010000101111011;  //       8571 
        86: sine = 18'b000010000111011110;  //       8670 
        87: sine = 18'b000010001001000010;  //       8770 
        88: sine = 18'b000010001010100110;  //       8870 
        89: sine = 18'b000010001100001001;  //       8969 
        90: sine = 18'b000010001101101101;  //       9069 
        91: sine = 18'b000010001111010000;  //       9168 
        92: sine = 18'b000010010000110100;  //       9268 
        93: sine = 18'b000010010010010111;  //       9367 
        94: sine = 18'b000010010011111011;  //       9467 
        95: sine = 18'b000010010101011110;  //       9566 
        96: sine = 18'b000010010111000010;  //       9666 
        97: sine = 18'b000010011000100101;  //       9765 
        98: sine = 18'b000010011010001001;  //       9865 
        99: sine = 18'b000010011011101100;  //       9964 
       100: sine = 18'b000010011101001111;  //      10063 
       101: sine = 18'b000010011110110011;  //      10163 
       102: sine = 18'b000010100000010110;  //      10262 
       103: sine = 18'b000010100001111001;  //      10361 
       104: sine = 18'b000010100011011101;  //      10461 
       105: sine = 18'b000010100101000000;  //      10560 
       106: sine = 18'b000010100110100011;  //      10659 
       107: sine = 18'b000010101000000110;  //      10758 
       108: sine = 18'b000010101001101001;  //      10857 
       109: sine = 18'b000010101011001100;  //      10956 
       110: sine = 18'b000010101100110000;  //      11056 
       111: sine = 18'b000010101110010011;  //      11155 
       112: sine = 18'b000010101111110110;  //      11254 
       113: sine = 18'b000010110001011001;  //      11353 
       114: sine = 18'b000010110010111100;  //      11452 
       115: sine = 18'b000010110100011111;  //      11551 
       116: sine = 18'b000010110110000010;  //      11650 
       117: sine = 18'b000010110111100101;  //      11749 
       118: sine = 18'b000010111001000111;  //      11847 
       119: sine = 18'b000010111010101010;  //      11946 
       120: sine = 18'b000010111100001101;  //      12045 
       121: sine = 18'b000010111101110000;  //      12144 
       122: sine = 18'b000010111111010011;  //      12243 
       123: sine = 18'b000011000000110101;  //      12341 
       124: sine = 18'b000011000010011000;  //      12440 
       125: sine = 18'b000011000011111011;  //      12539 
       126: sine = 18'b000011000101011110;  //      12638 
       127: sine = 18'b000011000111000000;  //      12736 
       128: sine = 18'b000011001000100011;  //      12835 
       129: sine = 18'b000011001010000101;  //      12933 
       130: sine = 18'b000011001011101000;  //      13032 
       131: sine = 18'b000011001101001010;  //      13130 
       132: sine = 18'b000011001110101101;  //      13229 
       133: sine = 18'b000011010000001111;  //      13327 
       134: sine = 18'b000011010001110010;  //      13426 
       135: sine = 18'b000011010011010100;  //      13524 
       136: sine = 18'b000011010100110110;  //      13622 
       137: sine = 18'b000011010110011001;  //      13721 
       138: sine = 18'b000011010111111011;  //      13819 
       139: sine = 18'b000011011001011101;  //      13917 
       140: sine = 18'b000011011011000000;  //      14016 
       141: sine = 18'b000011011100100010;  //      14114 
       142: sine = 18'b000011011110000100;  //      14212 
       143: sine = 18'b000011011111100110;  //      14310 
       144: sine = 18'b000011100001001000;  //      14408 
       145: sine = 18'b000011100010101010;  //      14506 
       146: sine = 18'b000011100100001100;  //      14604 
       147: sine = 18'b000011100101101110;  //      14702 
       148: sine = 18'b000011100111010000;  //      14800 
       149: sine = 18'b000011101000110010;  //      14898 
       150: sine = 18'b000011101010010100;  //      14996 
       151: sine = 18'b000011101011110110;  //      15094 
       152: sine = 18'b000011101101011000;  //      15192 
       153: sine = 18'b000011101110111001;  //      15289 
       154: sine = 18'b000011110000011011;  //      15387 
       155: sine = 18'b000011110001111101;  //      15485 
       156: sine = 18'b000011110011011110;  //      15582 
       157: sine = 18'b000011110101000000;  //      15680 
       158: sine = 18'b000011110110100010;  //      15778 
       159: sine = 18'b000011111000000011;  //      15875 
       160: sine = 18'b000011111001100101;  //      15973 
       161: sine = 18'b000011111011000110;  //      16070 
       162: sine = 18'b000011111100101000;  //      16168 
       163: sine = 18'b000011111110001001;  //      16265 
       164: sine = 18'b000011111111101010;  //      16362 
       165: sine = 18'b000100000001001100;  //      16460 
       166: sine = 18'b000100000010101101;  //      16557 
       167: sine = 18'b000100000100001110;  //      16654 
       168: sine = 18'b000100000101101111;  //      16751 
       169: sine = 18'b000100000111010001;  //      16849 
       170: sine = 18'b000100001000110010;  //      16946 
       171: sine = 18'b000100001010010011;  //      17043 
       172: sine = 18'b000100001011110100;  //      17140 
       173: sine = 18'b000100001101010101;  //      17237 
       174: sine = 18'b000100001110110110;  //      17334 
       175: sine = 18'b000100010000010111;  //      17431 
       176: sine = 18'b000100010001111000;  //      17528 
       177: sine = 18'b000100010011011001;  //      17625 
       178: sine = 18'b000100010100111001;  //      17721 
       179: sine = 18'b000100010110011010;  //      17818 
       180: sine = 18'b000100010111111011;  //      17915 
       181: sine = 18'b000100011001011100;  //      18012 
       182: sine = 18'b000100011010111100;  //      18108 
       183: sine = 18'b000100011100011101;  //      18205 
       184: sine = 18'b000100011101111101;  //      18301 
       185: sine = 18'b000100011111011110;  //      18398 
       186: sine = 18'b000100100000111110;  //      18494 
       187: sine = 18'b000100100010011111;  //      18591 
       188: sine = 18'b000100100011111111;  //      18687 
       189: sine = 18'b000100100101011111;  //      18783 
       190: sine = 18'b000100100111000000;  //      18880 
       191: sine = 18'b000100101000100000;  //      18976 
       192: sine = 18'b000100101010000000;  //      19072 
       193: sine = 18'b000100101011100000;  //      19168 
       194: sine = 18'b000100101101000000;  //      19264 
       195: sine = 18'b000100101110100001;  //      19361 
       196: sine = 18'b000100110000000001;  //      19457 
       197: sine = 18'b000100110001100001;  //      19553 
       198: sine = 18'b000100110011000000;  //      19648 
       199: sine = 18'b000100110100100000;  //      19744 
       200: sine = 18'b000100110110000000;  //      19840 
       201: sine = 18'b000100110111100000;  //      19936 
       202: sine = 18'b000100111001000000;  //      20032 
       203: sine = 18'b000100111010011111;  //      20127 
       204: sine = 18'b000100111011111111;  //      20223 
       205: sine = 18'b000100111101011111;  //      20319 
       206: sine = 18'b000100111110111110;  //      20414 
       207: sine = 18'b000101000000011110;  //      20510 
       208: sine = 18'b000101000001111101;  //      20605 
       209: sine = 18'b000101000011011101;  //      20701 
       210: sine = 18'b000101000100111100;  //      20796 
       211: sine = 18'b000101000110011011;  //      20891 
       212: sine = 18'b000101000111111011;  //      20987 
       213: sine = 18'b000101001001011010;  //      21082 
       214: sine = 18'b000101001010111001;  //      21177 
       215: sine = 18'b000101001100011000;  //      21272 
       216: sine = 18'b000101001101110111;  //      21367 
       217: sine = 18'b000101001111010110;  //      21462 
       218: sine = 18'b000101010000110101;  //      21557 
       219: sine = 18'b000101010010010100;  //      21652 
       220: sine = 18'b000101010011110011;  //      21747 
       221: sine = 18'b000101010101010010;  //      21842 
       222: sine = 18'b000101010110110000;  //      21936 
       223: sine = 18'b000101011000001111;  //      22031 
       224: sine = 18'b000101011001101110;  //      22126 
       225: sine = 18'b000101011011001100;  //      22220 
       226: sine = 18'b000101011100101011;  //      22315 
       227: sine = 18'b000101011110001001;  //      22409 
       228: sine = 18'b000101011111101000;  //      22504 
       229: sine = 18'b000101100001000110;  //      22598 
       230: sine = 18'b000101100010100101;  //      22693 
       231: sine = 18'b000101100100000011;  //      22787 
       232: sine = 18'b000101100101100001;  //      22881 
       233: sine = 18'b000101100110111111;  //      22975 
       234: sine = 18'b000101101000011101;  //      23069 
       235: sine = 18'b000101101001111011;  //      23163 
       236: sine = 18'b000101101011011001;  //      23257 
       237: sine = 18'b000101101100110111;  //      23351 
       238: sine = 18'b000101101110010101;  //      23445 
       239: sine = 18'b000101101111110011;  //      23539 
       240: sine = 18'b000101110001010001;  //      23633 
       241: sine = 18'b000101110010101111;  //      23727 
       242: sine = 18'b000101110100001100;  //      23820 
       243: sine = 18'b000101110101101010;  //      23914 
       244: sine = 18'b000101110111001000;  //      24008 
       245: sine = 18'b000101111000100101;  //      24101 
       246: sine = 18'b000101111010000011;  //      24195 
       247: sine = 18'b000101111011100000;  //      24288 
       248: sine = 18'b000101111100111101;  //      24381 
       249: sine = 18'b000101111110011011;  //      24475 
       250: sine = 18'b000101111111111000;  //      24568 
       251: sine = 18'b000110000001010101;  //      24661 
       252: sine = 18'b000110000010110010;  //      24754 
       253: sine = 18'b000110000100001111;  //      24847 
       254: sine = 18'b000110000101101100;  //      24940 
       255: sine = 18'b000110000111001001;  //      25033 
       256: sine = 18'b000110001000100110;  //      25126 
       257: sine = 18'b000110001010000011;  //      25219 
       258: sine = 18'b000110001011100000;  //      25312 
       259: sine = 18'b000110001100111100;  //      25404 
       260: sine = 18'b000110001110011001;  //      25497 
       261: sine = 18'b000110001111110101;  //      25589 
       262: sine = 18'b000110010001010010;  //      25682 
       263: sine = 18'b000110010010101110;  //      25774 
       264: sine = 18'b000110010100001011;  //      25867 
       265: sine = 18'b000110010101100111;  //      25959 
       266: sine = 18'b000110010111000011;  //      26051 
       267: sine = 18'b000110011000100000;  //      26144 
       268: sine = 18'b000110011001111100;  //      26236 
       269: sine = 18'b000110011011011000;  //      26328 
       270: sine = 18'b000110011100110100;  //      26420 
       271: sine = 18'b000110011110010000;  //      26512 
       272: sine = 18'b000110011111101100;  //      26604 
       273: sine = 18'b000110100001001000;  //      26696 
       274: sine = 18'b000110100010100011;  //      26787 
       275: sine = 18'b000110100011111111;  //      26879 
       276: sine = 18'b000110100101011011;  //      26971 
       277: sine = 18'b000110100110110110;  //      27062 
       278: sine = 18'b000110101000010010;  //      27154 
       279: sine = 18'b000110101001101101;  //      27245 
       280: sine = 18'b000110101011001001;  //      27337 
       281: sine = 18'b000110101100100100;  //      27428 
       282: sine = 18'b000110101101111111;  //      27519 
       283: sine = 18'b000110101111011011;  //      27611 
       284: sine = 18'b000110110000110110;  //      27702 
       285: sine = 18'b000110110010010001;  //      27793 
       286: sine = 18'b000110110011101100;  //      27884 
       287: sine = 18'b000110110101000111;  //      27975 
       288: sine = 18'b000110110110100010;  //      28066 
       289: sine = 18'b000110110111111100;  //      28156 
       290: sine = 18'b000110111001010111;  //      28247 
       291: sine = 18'b000110111010110010;  //      28338 
       292: sine = 18'b000110111100001101;  //      28429 
       293: sine = 18'b000110111101100111;  //      28519 
       294: sine = 18'b000110111111000010;  //      28610 
       295: sine = 18'b000111000000011100;  //      28700 
       296: sine = 18'b000111000001110110;  //      28790 
       297: sine = 18'b000111000011010001;  //      28881 
       298: sine = 18'b000111000100101011;  //      28971 
       299: sine = 18'b000111000110000101;  //      29061 
       300: sine = 18'b000111000111011111;  //      29151 
       301: sine = 18'b000111001000111001;  //      29241 
       302: sine = 18'b000111001010010011;  //      29331 
       303: sine = 18'b000111001011101101;  //      29421 
       304: sine = 18'b000111001101000111;  //      29511 
       305: sine = 18'b000111001110100000;  //      29600 
       306: sine = 18'b000111001111111010;  //      29690 
       307: sine = 18'b000111010001010100;  //      29780 
       308: sine = 18'b000111010010101101;  //      29869 
       309: sine = 18'b000111010100000111;  //      29959 
       310: sine = 18'b000111010101100000;  //      30048 
       311: sine = 18'b000111010110111001;  //      30137 
       312: sine = 18'b000111011000010010;  //      30226 
       313: sine = 18'b000111011001101100;  //      30316 
       314: sine = 18'b000111011011000101;  //      30405 
       315: sine = 18'b000111011100011110;  //      30494 
       316: sine = 18'b000111011101110111;  //      30583 
       317: sine = 18'b000111011111010000;  //      30672 
       318: sine = 18'b000111100000101000;  //      30760 
       319: sine = 18'b000111100010000001;  //      30849 
       320: sine = 18'b000111100011011010;  //      30938 
       321: sine = 18'b000111100100110010;  //      31026 
       322: sine = 18'b000111100110001011;  //      31115 
       323: sine = 18'b000111100111100011;  //      31203 
       324: sine = 18'b000111101000111100;  //      31292 
       325: sine = 18'b000111101010010100;  //      31380 
       326: sine = 18'b000111101011101100;  //      31468 
       327: sine = 18'b000111101101000100;  //      31556 
       328: sine = 18'b000111101110011100;  //      31644 
       329: sine = 18'b000111101111110100;  //      31732 
       330: sine = 18'b000111110001001100;  //      31820 
       331: sine = 18'b000111110010100100;  //      31908 
       332: sine = 18'b000111110011111100;  //      31996 
       333: sine = 18'b000111110101010100;  //      32084 
       334: sine = 18'b000111110110101011;  //      32171 
       335: sine = 18'b000111111000000011;  //      32259 
       336: sine = 18'b000111111001011010;  //      32346 
       337: sine = 18'b000111111010110010;  //      32434 
       338: sine = 18'b000111111100001001;  //      32521 
       339: sine = 18'b000111111101100000;  //      32608 
       340: sine = 18'b000111111110110111;  //      32695 
       341: sine = 18'b001000000000001111;  //      32783 
       342: sine = 18'b001000000001100110;  //      32870 
       343: sine = 18'b001000000010111100;  //      32956 
       344: sine = 18'b001000000100010011;  //      33043 
       345: sine = 18'b001000000101101010;  //      33130 
       346: sine = 18'b001000000111000001;  //      33217 
       347: sine = 18'b001000001000010111;  //      33303 
       348: sine = 18'b001000001001101110;  //      33390 
       349: sine = 18'b001000001011000100;  //      33476 
       350: sine = 18'b001000001100011011;  //      33563 
       351: sine = 18'b001000001101110001;  //      33649 
       352: sine = 18'b001000001111000111;  //      33735 
       353: sine = 18'b001000010000011101;  //      33821 
       354: sine = 18'b001000010001110100;  //      33908 
       355: sine = 18'b001000010011001010;  //      33994 
       356: sine = 18'b001000010100011111;  //      34079 
       357: sine = 18'b001000010101110101;  //      34165 
       358: sine = 18'b001000010111001011;  //      34251 
       359: sine = 18'b001000011000100001;  //      34337 
       360: sine = 18'b001000011001110110;  //      34422 
       361: sine = 18'b001000011011001100;  //      34508 
       362: sine = 18'b001000011100100001;  //      34593 
       363: sine = 18'b001000011101110111;  //      34679 
       364: sine = 18'b001000011111001100;  //      34764 
       365: sine = 18'b001000100000100001;  //      34849 
       366: sine = 18'b001000100001110110;  //      34934 
       367: sine = 18'b001000100011001011;  //      35019 
       368: sine = 18'b001000100100100000;  //      35104 
       369: sine = 18'b001000100101110101;  //      35189 
       370: sine = 18'b001000100111001010;  //      35274 
       371: sine = 18'b001000101000011110;  //      35358 
       372: sine = 18'b001000101001110011;  //      35443 
       373: sine = 18'b001000101011000111;  //      35527 
       374: sine = 18'b001000101100011100;  //      35612 
       375: sine = 18'b001000101101110000;  //      35696 
       376: sine = 18'b001000101111000101;  //      35781 
       377: sine = 18'b001000110000011001;  //      35865 
       378: sine = 18'b001000110001101101;  //      35949 
       379: sine = 18'b001000110011000001;  //      36033 
       380: sine = 18'b001000110100010101;  //      36117 
       381: sine = 18'b001000110101101001;  //      36201 
       382: sine = 18'b001000110110111100;  //      36284 
       383: sine = 18'b001000111000010000;  //      36368 
       384: sine = 18'b001000111001100100;  //      36452 
       385: sine = 18'b001000111010110111;  //      36535 
       386: sine = 18'b001000111100001011;  //      36619 
       387: sine = 18'b001000111101011110;  //      36702 
       388: sine = 18'b001000111110110001;  //      36785 
       389: sine = 18'b001001000000000100;  //      36868 
       390: sine = 18'b001001000001010111;  //      36951 
       391: sine = 18'b001001000010101010;  //      37034 
       392: sine = 18'b001001000011111101;  //      37117 
       393: sine = 18'b001001000101010000;  //      37200 
       394: sine = 18'b001001000110100011;  //      37283 
       395: sine = 18'b001001000111110101;  //      37365 
       396: sine = 18'b001001001001001000;  //      37448 
       397: sine = 18'b001001001010011010;  //      37530 
       398: sine = 18'b001001001011101101;  //      37613 
       399: sine = 18'b001001001100111111;  //      37695 
       400: sine = 18'b001001001110010001;  //      37777 
       401: sine = 18'b001001001111100011;  //      37859 
       402: sine = 18'b001001010000110101;  //      37941 
       403: sine = 18'b001001010010000111;  //      38023 
       404: sine = 18'b001001010011011001;  //      38105 
       405: sine = 18'b001001010100101011;  //      38187 
       406: sine = 18'b001001010101111101;  //      38269 
       407: sine = 18'b001001010111001110;  //      38350 
       408: sine = 18'b001001011000100000;  //      38432 
       409: sine = 18'b001001011001110001;  //      38513 
       410: sine = 18'b001001011011000010;  //      38594 
       411: sine = 18'b001001011100010011;  //      38675 
       412: sine = 18'b001001011101100101;  //      38757 
       413: sine = 18'b001001011110110110;  //      38838 
       414: sine = 18'b001001100000000111;  //      38919 
       415: sine = 18'b001001100001010111;  //      38999 
       416: sine = 18'b001001100010101000;  //      39080 
       417: sine = 18'b001001100011111001;  //      39161 
       418: sine = 18'b001001100101001001;  //      39241 
       419: sine = 18'b001001100110011010;  //      39322 
       420: sine = 18'b001001100111101010;  //      39402 
       421: sine = 18'b001001101000111010;  //      39482 
       422: sine = 18'b001001101010001011;  //      39563 
       423: sine = 18'b001001101011011011;  //      39643 
       424: sine = 18'b001001101100101011;  //      39723 
       425: sine = 18'b001001101101111011;  //      39803 
       426: sine = 18'b001001101111001010;  //      39882 
       427: sine = 18'b001001110000011010;  //      39962 
       428: sine = 18'b001001110001101010;  //      40042 
       429: sine = 18'b001001110010111001;  //      40121 
       430: sine = 18'b001001110100001001;  //      40201 
       431: sine = 18'b001001110101011000;  //      40280 
       432: sine = 18'b001001110110100111;  //      40359 
       433: sine = 18'b001001110111110111;  //      40439 
       434: sine = 18'b001001111001000110;  //      40518 
       435: sine = 18'b001001111010010101;  //      40597 
       436: sine = 18'b001001111011100011;  //      40675 
       437: sine = 18'b001001111100110010;  //      40754 
       438: sine = 18'b001001111110000001;  //      40833 
       439: sine = 18'b001001111111010000;  //      40912 
       440: sine = 18'b001010000000011110;  //      40990 
       441: sine = 18'b001010000001101100;  //      41068 
       442: sine = 18'b001010000010111011;  //      41147 
       443: sine = 18'b001010000100001001;  //      41225 
       444: sine = 18'b001010000101010111;  //      41303 
       445: sine = 18'b001010000110100101;  //      41381 
       446: sine = 18'b001010000111110011;  //      41459 
       447: sine = 18'b001010001001000001;  //      41537 
       448: sine = 18'b001010001010001110;  //      41614 
       449: sine = 18'b001010001011011100;  //      41692 
       450: sine = 18'b001010001100101010;  //      41770 
       451: sine = 18'b001010001101110111;  //      41847 
       452: sine = 18'b001010001111000100;  //      41924 
       453: sine = 18'b001010010000010010;  //      42002 
       454: sine = 18'b001010010001011111;  //      42079 
       455: sine = 18'b001010010010101100;  //      42156 
       456: sine = 18'b001010010011111001;  //      42233 
       457: sine = 18'b001010010101000101;  //      42309 
       458: sine = 18'b001010010110010010;  //      42386 
       459: sine = 18'b001010010111011111;  //      42463 
       460: sine = 18'b001010011000101011;  //      42539 
       461: sine = 18'b001010011001111000;  //      42616 
       462: sine = 18'b001010011011000100;  //      42692 
       463: sine = 18'b001010011100010000;  //      42768 
       464: sine = 18'b001010011101011100;  //      42844 
       465: sine = 18'b001010011110101000;  //      42920 
       466: sine = 18'b001010011111110100;  //      42996 
       467: sine = 18'b001010100001000000;  //      43072 
       468: sine = 18'b001010100010001100;  //      43148 
       469: sine = 18'b001010100011010111;  //      43223 
       470: sine = 18'b001010100100100011;  //      43299 
       471: sine = 18'b001010100101101110;  //      43374 
       472: sine = 18'b001010100110111010;  //      43450 
       473: sine = 18'b001010101000000101;  //      43525 
       474: sine = 18'b001010101001010000;  //      43600 
       475: sine = 18'b001010101010011011;  //      43675 
       476: sine = 18'b001010101011100110;  //      43750 
       477: sine = 18'b001010101100110001;  //      43825 
       478: sine = 18'b001010101101111011;  //      43899 
       479: sine = 18'b001010101111000110;  //      43974 
       480: sine = 18'b001010110000010001;  //      44049 
       481: sine = 18'b001010110001011011;  //      44123 
       482: sine = 18'b001010110010100101;  //      44197 
       483: sine = 18'b001010110011101111;  //      44271 
       484: sine = 18'b001010110100111001;  //      44345 
       485: sine = 18'b001010110110000011;  //      44419 
       486: sine = 18'b001010110111001101;  //      44493 
       487: sine = 18'b001010111000010111;  //      44567 
       488: sine = 18'b001010111001100001;  //      44641 
       489: sine = 18'b001010111010101010;  //      44714 
       490: sine = 18'b001010111011110100;  //      44788 
       491: sine = 18'b001010111100111101;  //      44861 
       492: sine = 18'b001010111110000110;  //      44934 
       493: sine = 18'b001010111111001111;  //      45007 
       494: sine = 18'b001011000000011000;  //      45080 
       495: sine = 18'b001011000001100001;  //      45153 
       496: sine = 18'b001011000010101010;  //      45226 
       497: sine = 18'b001011000011110011;  //      45299 
       498: sine = 18'b001011000100111011;  //      45371 
       499: sine = 18'b001011000110000100;  //      45444 
       500: sine = 18'b001011000111001100;  //      45516 
       501: sine = 18'b001011001000010101;  //      45589 
       502: sine = 18'b001011001001011101;  //      45661 
       503: sine = 18'b001011001010100101;  //      45733 
       504: sine = 18'b001011001011101101;  //      45805 
       505: sine = 18'b001011001100110101;  //      45877 
       506: sine = 18'b001011001101111100;  //      45948 
       507: sine = 18'b001011001111000100;  //      46020 
       508: sine = 18'b001011010000001011;  //      46091 
       509: sine = 18'b001011010001010011;  //      46163 
       510: sine = 18'b001011010010011010;  //      46234 
       511: sine = 18'b001011010011100001;  //      46305 
    endcase 
endmodule 


