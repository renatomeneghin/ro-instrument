// -----------------------------------------------------------------------------
//Actel Corporation Proprietary and Confidential
//Copyright 2008 Actel Corporation. All rights reserved.
//
//ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
//ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
//IN ADVANCE IN WRITING.
//
//Description:  CoreFFT RTL 
//              Customized Twiddle Coefficients 
//
//Revision Information:
//Date         Description
//05Nov2009    Initial Release 
//
//SVN Revision Information:
//SVN $Revision: $
//SVN $Data: $
//
//Resolved SARs
//SAR     Date    Who         Description
//
//Notes:

`timescale 1 ns/100 ps

module COREFFT_C1_COREFFT_C1_0_twiddle (A,T);
  parameter TDWIDTH = 16;
  parameter LOGPTS  = 5;

  input	[LOGPTS-2:0]	A;	// Address
  output reg [TDWIDTH-1:0]	T;	// Table output

  always @ (A)
    case (A) // synopsys parallel_case
      9'h0: T=64'b0000000000000000000000000000000001111111111111111111111111111111;  //     0 2147483647
      9'h1: T=64'b0000000011001001000011111000100001111111111111110110001000010101;  // 13176712 2147443221
      9'h2: T=64'b0000000110010010000111010010000001111111111111011000100001011001;  // 26352928 2147321945
      9'h3: T=64'b0000001001011011001001101101011101111111111110100111001011010000;  // 39528151 2147119824
      9'h4: T=64'b0000001100100100001010101011111101111111111101100010000110000001;  // 52701887 2146836865
      9'h5: T=64'b0000001111101101001001101110011001111111111100001001010001110111;  // 65873638 2146473079
      9'h6: T=64'b0000010010110110000110010101110101111111111010011100101110111111;  // 79042909 2146028479
      9'h7: T=64'b0000010101111111000000000011010101111111111000011100011101101010;  // 92209205 2145503082
      9'h8: T=64'b0000011001000111110110010111110001111111110110001000011110001101;  // 105372028 2144896909
      9'h9: T=64'b0000011100010000101000110100010101111111110011100000110000111101;  // 118530885 2144209981
      9'ha: T=64'b0000011111011001010110111001111001111111110000100101010110010101;  // 131685278 2143442325
      9'hb: T=64'b0000100010100010000000001001101001111111101101010110001110110010;  // 144834714 2142593970
      9'hc: T=64'b0000100101101010100100000100100101111111101001110011011010110011;  // 157978697 2141664947
      9'hd: T=64'b0000101000110011000010001011110001111111100101111100111010111100;  // 171116732 2140655292
      9'he: T=64'b0000101011111011011010000000010101111111100001110010101111110010;  // 184248325 2139565042
      9'hf: T=64'b0000101111000011101011000011010101111111011101010100111001111111;  // 197372981 2138394239
      9'h10: T=64'b0000110010001011110100110101111001111111011000100011011010001110;  // 210490206 2137142926
      9'h11: T=64'b0000110101010011110110111001001001111111010011011110010001010000;  // 223599506 2135811152
      9'h12: T=64'b0000111000011011110000101110010001111111001110000101011111110101;  // 236700388 2134398965
      9'h13: T=64'b0000111011100011100001110110011001111111001000011001000110110011;  // 249792358 2132906419
      9'h14: T=64'b0000111110101011001001110010101101111111000010011001000111000011;  // 262874923 2131333571
      9'h15: T=64'b0001000001110010101000000100100001111110111100000101100001011111;  // 275947592 2129680479
      9'h16: T=64'b0001000100111001111100001100111101111110110101011110010111000101;  // 289009871 2127947205
      9'h17: T=64'b0001001000000001000101101101010101111110101110100011101000111000;  // 302061269 2126133816
      9'h18: T=64'b0001001011001000000100000110111001111110100111010101010111111011;  // 315101294 2124240379
      9'h19: T=64'b0001001110001110110110111011000101111110011111110011100101010110;  // 328129457 2122266966
      9'h1a: T=64'b0001010001010101011101101011000101111110010111111110010010010010;  // 341145265 2120213650
      9'h1b: T=64'b0001010100011011110111111000010101111110001111110101011111111110;  // 354148229 2118080510
      9'h1c: T=64'b0001010111100010000101000100010001111110000111011001001111101001;  // 367137860 2115867625
      9'h1d: T=64'b0001011010101000000100110000010101111101111110101001100010100111;  // 380113669 2113575079
      9'h1e: T=64'b0001011101101101110110011101111001111101110101100110011010001110;  // 393075166 2111202958
      9'h1f: T=64'b0001100000110011011001101110100001111101101100001111110111110111;  // 406021864 2108751351
      9'h20: T=64'b0001100011111000101110000011110001111101100010100101111100111111;  // 418953276 2106220351
      9'h21: T=64'b0001100110111101110010111111001101111101011000101000101011000101;  // 431868915 2103610053
      9'h22: T=64'b0001101010000010101000000010010101111101001110011000000011101011;  // 444768293 2100920555
      9'h23: T=64'b0001101101000111001100101110111101111101000011110100001000010111;  // 457650927 2098151959
      9'h24: T=64'b0001110000001011100000100110101001111100111000111100111010110001;  // 470516330 2095304369
      9'h25: T=64'b0001110011001111100011001011001101111100101101110010011100100011;  // 483364019 2092377891
      9'h26: T=64'b0001110110010011010011111110010101111100100010010100101111011101;  // 496193509 2089372637
      9'h27: T=64'b0001111001010110110010100001111001111100010110100011110101001111;  // 509004318 2086288719
      9'h28: T=64'b0001111100011001111110010111101101111100001010011111101111101101;  // 521795963 2083126253
      9'h29: T=64'b0001111111011100110111000001101101111011111110001000100000101111;  // 534567963 2079885359
      9'h2a: T=64'b0010000010011111011100000001110001111011110001011110001010001111;  // 547319836 2076566159
      9'h2b: T=64'b0010000101100001101100111001111101111011100100100000101110001000;  // 560051103 2073168776
      9'h2c: T=64'b0010001000100011101001001100010101111011010111010000001110011101;  // 572761285 2069693341
      9'h2d: T=64'b0010001011100101010000011010111101111011001001101100101101001110;  // 585449903 2066139982
      9'h2e: T=64'b0010001110100110100010000111111001111010111011110110001100100011;  // 598116478 2062508835
      9'h2f: T=64'b0010010001100111011101110101011101111010101101101100101110100011;  // 610760535 2058800035
      9'h30: T=64'b0010010100101000000011000101110101111010011111010000010101011010;  // 623381597 2055013722
      9'h31: T=64'b0010010111101000010001011011011001111010010000100001000011011000;  // 635979190 2051150040
      9'h32: T=64'b0010011010101000001000011000010101111010000001011110111010101100;  // 648552837 2047209132
      9'h33: T=64'b0010011101100111100111011111010001111001110010001001111101101101;  // 661102068 2043191149
      9'h34: T=64'b0010100000100110101110010010100001111001100010100010001110110000;  // 673626408 2039096240
      9'h35: T=64'b0010100011100101011100010100101001111001010010100111110000010001;  // 686125386 2034924561
      9'h36: T=64'b0010100110100011110001001000010101111001000010011010100100101100;  // 698598533 2030676268
      9'h37: T=64'b0010101001100001101100010000000101111000110001111010101110100001;  // 711045377 2026351521
      9'h38: T=64'b0010101100011111001101001110101101111000100001001000010000010011;  // 723465451 2021950483
      9'h39: T=64'b0010101111011100010011100110111101111000010000000011001100101000;  // 735858287 2017473320
      9'h3a: T=64'b0010110010011000111110111011101001110111111110101011100110001000;  // 748223418 2012920200
      9'h3b: T=64'b0010110101010101001110101111101101110111101101000001011111011111;  // 760560379 2008291295
      9'h3c: T=64'b0010111000010001000010100110001001110111011011000100111011011010;  // 772868706 2003586778
      9'h3d: T=64'b0010111011001100011010000001111001110111001000110101111100101100;  // 785147934 1998806828
      9'h3e: T=64'b0010111110000111010100100110001001110110110110010100100110001000;  // 797397602 1993951624
      9'h3f: T=64'b0011000001000001110001110110000001110110100011100000111010100101;  // 809617248 1989021349
      9'h40: T=64'b0011000011111011110001010100110101110110010000011010111100111100;  // 821806413 1984016188
      9'h41: T=64'b0011000110110101010010100101110101110101111101000010110000001010;  // 833964637 1978936330
      9'h42: T=64'b0011001001101110010101001100011101110101101001011000010111001110;  // 846091463 1973781966
      9'h43: T=64'b0011001100100110111000101100001001110101010101011011110101001011;  // 858186434 1968553291
      9'h44: T=64'b0011001111011110111100101000011101110101000001001101001101000100;  // 870249095 1963250500
      9'h45: T=64'b0011010010010110100000100100111101110100101100101100100010000011;  // 882278991 1957873795
      9'h46: T=64'b0011010101001101100100000101011001110100010111111001110111010000;  // 894275670 1952423376
      9'h47: T=64'b0011011000000100000110101101100101110100000010110101001111111010;  // 906238681 1946899450
      9'h48: T=64'b0011011010111010001000000001001101110011101101011110101111010000;  // 918167571 1941302224
      9'h49: T=64'b0011011101101111100111100100011001110011010111110110011000100101;  // 930061894 1935631909
      9'h4a: T=64'b0011100000100100100100111011000001110011000001111100001111001111;  // 941921200 1929888719
      9'h4b: T=64'b0011100011011000111111101001001101110010101011110000010110100110;  // 953745043 1924072870
      9'h4c: T=64'b0011100110001100110111010011001001110010010101010010110010000100;  // 965532978 1918184580
      9'h4d: T=64'b0011101001000000001011011101000101110001111110100011100101001000;  // 977284561 1912224072
      9'h4e: T=64'b0011101011110010111011101011011101110001100111100010110011010001;  // 988999351 1906191569
      9'h4f: T=64'b0011101110100101000111100010100101110001010000010000100000000100;  // 1000676905 1900087300
      9'h50: T=64'b0011110001010110101110100111000001110000111000101100101111000101;  // 1012316784 1893911493
      9'h51: T=64'b0011110100000111110000011101010101110000100000110111100011111110;  // 1023918549 1887664382
      9'h52: T=64'b0011110110111000001100101010010101110000001000110001000010011001;  // 1035481765 1881346201
      9'h53: T=64'b0011111001101000000010110010110001101111110000011001001110000100;  // 1047005996 1874957188
      9'h54: T=64'b0011111100010111010010011011011101101111010111110000001010110001;  // 1058490807 1868497585
      9'h55: T=64'b0011111111000101111011001001011101101110111110110101111100010001;  // 1069935767 1861967633
      9'h56: T=64'b0100000001110011111100100001110101101110100101101010100110011100;  // 1081340445 1855367580
      9'h57: T=64'b0100000100100001010110001001101001101110001100001110001101001001;  // 1092704410 1848697673
      9'h58: T=64'b0100000111001110000111100110010001101101110010100000110100010100;  // 1104027236 1841958164
      9'h59: T=64'b0100001001111010010000011101000001101101011000100010011111111001;  // 1115308496 1835149305
      9'h5a: T=64'b0100001100100101110000010011010101101100111110010011010011111011;  // 1126547765 1828271355
      9'h5b: T=64'b0100001111010000100110101110110001101100100011110011010100011011;  // 1137744620 1821324571
      9'h5c: T=64'b0100010001111010110011010101000001101100001001000010100101011111;  // 1148898640 1814309215
      9'h5d: T=64'b0100010100100100010101101011110001101011101110000001001011010000;  // 1160009404 1807225552
      9'h5e: T=64'b0100010111001101001101011000111101101011010010101111001001111000;  // 1171076495 1800073848
      9'h5f: T=64'b0100011001110101011010000010011101101010110111001100100101100100;  // 1182099495 1792854372
      9'h60: T=64'b0100011100011100111011001110011001101010011011011001100010100011;  // 1193077990 1785567395
      9'h61: T=64'b0100011111000011110000100010111001101001111111010110000101001010;  // 1204011566 1778213194
      9'h62: T=64'b0100100001101001111001100110010001101001100011000010010001101011;  // 1214899812 1770792043
      9'h63: T=64'b0100100100001111010101111110111001101001000110011110001100011111;  // 1225742318 1763304223
      9'h64: T=64'b0100100110110100000101010011001101101000101001101001111010000000;  // 1236538675 1755750016
      9'h65: T=64'b0100101001011000000111001001110101101000001100100101011110101010;  // 1247288477 1748129706
      9'h66: T=64'b0100101011111011011011001001011101100111101111010000111110111100;  // 1257991319 1740443580
      9'h67: T=64'b0100101110011110000000111000111101100111010001101100011111010111;  // 1268646799 1732691927
      9'h68: T=64'b0100110000111111110111111111001101100110110011111000000100011111;  // 1279254515 1724875039
      9'h69: T=64'b0100110011100001000000000011010001100110010101110011110010111011;  // 1289814068 1716993211
      9'h6a: T=64'b0100110110000001011000101100001101100101110111011111101111010010;  // 1300325059 1709046738
      9'h6b: T=64'b0100111000100001000001100001011101100101011000111011111110010001;  // 1310787095 1701035921
      9'h6c: T=64'b0100111010111111111010001010010001100100111010001000100100100101;  // 1321199780 1692961061
      9'h6d: T=64'b0100111101011110000010001110001001100100011011000101100110111111;  // 1331562722 1684822463
      9'h6e: T=64'b0100111111111011011001010100110001100011111011110011001010001111;  // 1341875532 1676620431
      9'h6f: T=64'b0101000010010111111111000101111001100011011100010001010011001100;  // 1352137822 1668355276
      9'h70: T=64'b0101000100110011110011001001010001100010111100100000000110101100;  // 1362349204 1660027308
      9'h71: T=64'b0101000111001110110101000110111001100010011100011111101001101000;  // 1372509294 1651636840
      9'h72: T=64'b0101001001101001000100100110111001100001111100010000000000111110;  // 1382617710 1643184190
      9'h73: T=64'b0101001100000010100001010001011101100001011011110001010001101011;  // 1392674071 1634669675
      9'h74: T=64'b0101001110011011001010101110111101100000111011000011100000101111;  // 1402677999 1626093615
      9'h75: T=64'b0101010000110011000000100111110101100000011010000110110011001110;  // 1412629117 1617456334
      9'h76: T=64'b0101010011001010000010100100101001011111111000111011001110001101;  // 1422527050 1608758157
      9'h77: T=64'b0101010101100000010000001110001001011111010111100000110110110010;  // 1432371426 1599999410
      9'h78: T=64'b0101010111110101101001001101001001011110110101110111110010001001;  // 1442161874 1591180425
      9'h79: T=64'b0101011010001010001101001010100101011110010100000000000101011101;  // 1451898025 1582301533
      9'h7a: T=64'b0101011100011101111011101111100101011101110001111001110101111011;  // 1461579513 1573363067
      9'h7b: T=64'b0101011110110000110100100101010101011101001111100101001000110110;  // 1471205973 1564365366
      9'h7c: T=64'b0101100001000010110111010101010001011100101101000010000011011111;  // 1480777044 1555308767
      9'h7d: T=64'b0101100011010100000011101000110001011100001010010000101011001100;  // 1490292364 1546193612
      9'h7e: T=64'b0101100101100100011001001001011101011011100111010001000101010011;  // 1499751575 1537020243
      9'h7f: T=64'b0101100111110011110111100001001001011011000100000011010111001110;  // 1509154322 1527789006
      9'h80: T=64'b0101101010000010011110011001100101011010100000100111100110011001;  // 1518500249 1518500249
      9'h81: T=64'b0101101100010000001101011100111001011001111100111101111000010010;  // 1527789006 1509154322
      9'h82: T=64'b0101101110011101000100010101001101011001011001000110010010010111;  // 1537020243 1499751575
      9'h83: T=64'b0101110000101001000010101100110001011000110101000000111010001100;  // 1546193612 1490292364
      9'h84: T=64'b0101110010110100001000001101111101011000010000101101110101010100;  // 1555308767 1480777044
      9'h85: T=64'b0101110100111110010100100011011001010111101100001101001001010101;  // 1564365366 1471205973
      9'h86: T=64'b0101110111000111100111010111101101010111000111011110111011111001;  // 1573363067 1461579513
      9'h87: T=64'b0101111001010000000000010101110101010110100010100011010010101001;  // 1582301533 1451898025
      9'h88: T=64'b0101111011010111011111001000100101010101111101011010010011010010;  // 1591180425 1442161874
      9'h89: T=64'b0101111101011110000011011011001001010101011000000100000011100010;  // 1599999410 1432371426
      9'h8a: T=64'b0101111111100011101100111000110101010100110010100000101001001010;  // 1608758157 1422527050
      9'h8b: T=64'b0110000001101000011011001100111001010100001100110000001001111101;  // 1617456334 1412629117
      9'h8c: T=64'b0110000011101100001110000010111101010011100110110010101011101111;  // 1626093615 1402677999
      9'h8d: T=64'b0110000101101111000101000110101101010011000000101000010100010111;  // 1634669675 1392674071
      9'h8e: T=64'b0110000111110001000000000011111001010010011010010001001001101110;  // 1643184190 1382617710
      9'h8f: T=64'b0110001001110001111110100110100001010001110011101101010001101110;  // 1651636840 1372509294
      9'h90: T=64'b0110001011110010000000011010110001010001001100111100110010010100;  // 1660027308 1362349204
      9'h91: T=64'b0110001101110001000101001100110001010000100101111111110001011110;  // 1668355276 1352137822
      9'h92: T=64'b0110001111101111001100101000111101001111111110110110010101001100;  // 1676620431 1341875532
      9'h93: T=64'b0110010001101100010110011011111101001111010111100000100011100010;  // 1684822463 1331562722
      9'h94: T=64'b0110010011101000100010010010010101001110101111111110100010100100;  // 1692961061 1321199780
      9'h95: T=64'b0110010101100011101111111001000101001110001000010000011000010111;  // 1701035921 1310787095
      9'h96: T=64'b0110010111011101111110111101001001001101100000010110001011000011;  // 1709046738 1300325059
      9'h97: T=64'b0110011001010111001111001011101101001100111000010000000000110100;  // 1716993211 1289814068
      9'h98: T=64'b0110011011001111100000010001111101001100001111111101111111110011;  // 1724875039 1279254515
      9'h99: T=64'b0110011101000110110001111101011101001011100111100000001110001111;  // 1732691927 1268646799
      9'h9a: T=64'b0110011110111101000011111011110001001010111110110110110010010111;  // 1740443580 1257991319
      9'h9b: T=64'b0110100000110010010101111010101001001010010110000001110010011101;  // 1748129706 1247288477
      9'h9c: T=64'b0110100010100110100111101000000001001001101101000001010100110011;  // 1755750016 1236538675
      9'h9d: T=64'b0110100100011001111000110001111101001001000011110101011111101110;  // 1763304223 1225742318
      9'h9e: T=64'b0110100110001100001001000110101101001000011010011110011001100100;  // 1770792043 1214899812
      9'h9f: T=64'b0110100111111101011000010100101001000111110000111100001000101110;  // 1778213194 1204011566
      9'ha0: T=64'b0110101001101101100110001010001101000111000111001110110011100110;  // 1785567395 1193077990
      9'ha1: T=64'b0110101011011100110010010110010001000110011101010110100000100111;  // 1792854372 1182099495
      9'ha2: T=64'b0110101101001010111100100111100001000101110011010011010110001111;  // 1800073848 1171076495
      9'ha3: T=64'b0110101110111000000100101101000001000101001001000101011010111100;  // 1807225552 1160009404
      9'ha4: T=64'b0110110000100100001010010101111101000100011110101100110101010000;  // 1814309215 1148898640
      9'ha5: T=64'b0110110010001111001101010001101101000011110100001001101011101100;  // 1821324571 1137744620
      9'ha6: T=64'b0110110011111001001101001111101101000011001001011100000100110101;  // 1828271355 1126547765
      9'ha7: T=64'b0110110101100010001001111111100101000010011110100100000111010000;  // 1835149305 1115308496
      9'ha8: T=64'b0110110111001010000011010001010001000001110011100001111001100100;  // 1841958164 1104027236
      9'ha9: T=64'b0110111000110000111000110100100101000001001000010101100010011010;  // 1848697673 1092704410
      9'haa: T=64'b0110111010010110101010011001110001000000011100111111001000011101;  // 1855367580 1081340445
      9'hab: T=64'b0110111011111011010111110001000100111111110001011110110010010111;  // 1861967633 1069935767
      9'hac: T=64'b0110111101011111000000101011000100111111000101110100100110110111;  // 1868497585 1058490807
      9'had: T=64'b0110111111000001100100111000010000111110011010000000101100101100;  // 1874957188 1047005996
      9'hae: T=64'b0111000000100011000100001001100100111101101110000011001010100101;  // 1881346201 1035481765
      9'haf: T=64'b0111000010000011011110001111111000111101000001111100000111010101;  // 1887664382 1023918549
      9'hb0: T=64'b0111000011100010110010111100010100111100010101101011101001110000;  // 1893911493 1012316784
      9'hb1: T=64'b0111000101000001000010000000010000111011101001010001111000101001;  // 1900087300 1000676905
      9'hb2: T=64'b0111000110011110001011001101000100111010111100101110111010110111;  // 1906191569 988999351
      9'hb3: T=64'b0111000111111010001110010100100000111010010000000010110111010001;  // 1912224072 977284561
      9'hb4: T=64'b0111001001010101001011001000010000111001100011001101110100110010;  // 1918184580 965532978
      9'hb5: T=64'b0111001010101111000001011010011000111000110110001111111010010011;  // 1924072870 953745043
      9'hb6: T=64'b0111001100000111110000111100111100111000001001001001001110110000;  // 1929888719 941921200
      9'hb7: T=64'b0111001101011111011001100010010100110111011011111001111001000110;  // 1935631909 930061894
      9'hb8: T=64'b0111001110110101111010111101000000110110101110100010000000010011;  // 1941302224 918167571
      9'hb9: T=64'b0111010000001011010100111111101000110110000001000001101011011001;  // 1946899450 906238681
      9'hba: T=64'b0111010001011111100111011101000000110101010011011001000001010110;  // 1952423376 894275670
      9'hbb: T=64'b0111010010110010110010001000001100110100100101101000001001001111;  // 1957873795 882278991
      9'hbc: T=64'b0111010100000100110100110100010000110011110111101111001010000111;  // 1963250500 870249095
      9'hbd: T=64'b0111010101010101101111010100101100110011001001101110001011000010;  // 1968553291 858186434
      9'hbe: T=64'b0111010110100101100001011100111000110010011011100101010011000111;  // 1973781966 846091463
      9'hbf: T=64'b0111010111110100001011000000101000110001101101010100101001011101;  // 1978936330 833964637
      9'hc0: T=64'b0111011001000001101011110011110000110000111110111100010101001101;  // 1984016188 821806413
      9'hc1: T=64'b0111011010001110000011101010010100110000010000011100011101100000;  // 1989021349 809617248
      9'hc2: T=64'b0111011011011001010010011000100000101111100001110101001001100010;  // 1993951624 797397602
      9'hc3: T=64'b0111011100100011010111110010110000101110110011000110100000011110;  // 1998806828 785147934
      9'hc4: T=64'b0111011101101100010011101101101000101110000100010000101001100010;  // 2003586778 772868706
      9'hc5: T=64'b0111011110110100000101111101111100101101010101010011101011111011;  // 2008291295 760560379
      9'hc6: T=64'b0111011111111010101110011000100000101100100110001111101110111010;  // 2012920200 748223418
      9'hc7: T=64'b0111100001000000001100110010100000101011110111000100111001101111;  // 2017473320 735858287
      9'hc8: T=64'b0111100010000100100001000001001100101011000111110011010011101011;  // 2021950483 723465451
      9'hc9: T=64'b0111100011000111101010111010000100101010011000011011000100000001;  // 2026351521 711045377
      9'hca: T=64'b0111100100001001101010010010110000101001101000111100010010000101;  // 2030676268 698598533
      9'hcb: T=64'b0111100101001010011111000001000100101000111001010111000101001010;  // 2034924561 686125386
      9'hcc: T=64'b0111100110001010001000111011000000101000001001101011100100101000;  // 2039096240 673626408
      9'hcd: T=64'b0111100111001000100111110110110100100111011001111001110111110100;  // 2043191149 661102068
      9'hce: T=64'b0111101000000101111011101010110000100110101010000010000110000101;  // 2047209132 648552837
      9'hcf: T=64'b0111101001000010000100001101100000100101111010000100010110110110;  // 2051150040 635979190
      9'hd0: T=64'b0111101001111101000001010101101000100101001010000000110001011101;  // 2055013722 623381597
      9'hd1: T=64'b0111101010110110110010111010001100100100011001110111011101010111;  // 2058800035 610760535
      9'hd2: T=64'b0111101011101111011000110010001100100011101001101000100001111110;  // 2062508835 598116478
      9'hd3: T=64'b0111101100100110110010110100111000100010111001010100000110101111;  // 2066139982 585449903
      9'hd4: T=64'b0111101101011101000000111001110100100010001000111010010011000101;  // 2069693341 572761285
      9'hd5: T=64'b0111101110010010000010111000100000100001011000011011001110011111;  // 2073168776 560051103
      9'hd6: T=64'b0111101111000101111000101000111100100000100111110111000000011100;  // 2076566159 547319836
      9'hd7: T=64'b0111101111111000100010000010111100011111110111001101110000011011;  // 2079885359 534567963
      9'hd8: T=64'b0111110000101001111110111110110100011111000110011111100101111011;  // 2083126253 521795963
      9'hd9: T=64'b0111110001011010001111010100111100011110010101101100101000011110;  // 2086288719 509004318
      9'hda: T=64'b0111110010001001010010111101110100011101100100110100111111100101;  // 2089372637 496193509
      9'hdb: T=64'b0111110010110111001001110010001100011100110011111000110010110011;  // 2092377891 483364019
      9'hdc: T=64'b0111110011100011110011101011000100011100000010111000001001101010;  // 2095304369 470516330
      9'hdd: T=64'b0111110100001111010000100001011100011011010001110011001011101111;  // 2098151959 457650927
      9'hde: T=64'b0111110100111001100000001110101100011010100000101010000000100101;  // 2100920555 444768293
      9'hdf: T=64'b0111110101100010100010101100010100011001101111011100101111110011;  // 2103610053 431868915
      9'he0: T=64'b0111110110001010010111110011111100011000111110001011100000111100;  // 2106220351 418953276
      9'he1: T=64'b0111110110110000111111011111011100011000001100110110011011101000;  // 2108751351 406021864
      9'he2: T=64'b0111110111010110011001101000111000010111011011011101100111011110;  // 2111202958 393075166
      9'he3: T=64'b0111110111111010100110001010011100010110101010000001001100000101;  // 2113575079 380113669
      9'he4: T=64'b0111111000011101100100111110100100010101111000100001010001000100;  // 2115867625 367137860
      9'he5: T=64'b0111111000111111010101111111111000010101000110111101111110000101;  // 2118080510 354148229
      9'he6: T=64'b0111111001011111111001001001001000010100010101010111011010110001;  // 2120213650 341145265
      9'he7: T=64'b0111111001111111001110010101011000010011100011101101101110110001;  // 2122266966 328129457
      9'he8: T=64'b0111111010011101010101011111101100010010110010000001000001101110;  // 2124240379 315101294
      9'he9: T=64'b0111111010111010001110100011100000010010000000010001011011010101;  // 2126133816 302061269
      9'hea: T=64'b0111111011010101111001011100010100010001001110011111000011001111;  // 2127947205 289009871
      9'heb: T=64'b0111111011110000010110000101111100010000011100101010000001001000;  // 2129680479 275947592
      9'hec: T=64'b0111111100001001100100011100001100001111101010110010011100101011;  // 2131333571 262874923
      9'hed: T=64'b0111111100100001100100011011001100001110111000111000011101100110;  // 2132906419 249792358
      9'hee: T=64'b0111111100111000010101111111010100001110000110111100001011100100;  // 2134398965 236700388
      9'hef: T=64'b0111111101001101111001000101000000001101010100111101101110010010;  // 2135811152 223599506
      9'hf0: T=64'b0111111101100010001101101000111000001100100010111101001101011110;  // 2137142926 210490206
      9'hf1: T=64'b0111111101110101010011100111111100001011110000111010110000110101;  // 2138394239 197372981
      9'hf2: T=64'b0111111110000111001010111111001000001010111110110110100000000101;  // 2139565042 184248325
      9'hf3: T=64'b0111111110010111110011101011110000001010001100110000100010111100;  // 2140655292 171116732
      9'hf4: T=64'b0111111110100111001101101011001100001001011010101001000001001001;  // 2141664947 157978697
      9'hf5: T=64'b0111111110110101011000111011001000001000101000100000000010011010;  // 2142593970 144834714
      9'hf6: T=64'b0111111111000010010101011001010100000111110110010101101110011110;  // 2143442325 131685278
      9'hf7: T=64'b0111111111001110000011000011110100000111000100001010001101000101;  // 2144209981 118530885
      9'hf8: T=64'b0111111111011000100001111000110100000110010001111101100101111100;  // 2144896909 105372028
      9'hf9: T=64'b0111111111100001110001110110101000000101011111110000000000110101;  // 2145503082 92209205
      9'hfa: T=64'b0111111111101001110010111011111100000100101101100001100101011101;  // 2146028479 79042909
      9'hfb: T=64'b0111111111110000100101000111011100000011111011010010011011100110;  // 2146473079 65873638
      9'hfc: T=64'b0111111111110110001000011000000100000011001001000010101010111111;  // 2146836865 52701887
      9'hfd: T=64'b0111111111111010011100101101000000000010010110110010011011010111;  // 2147119824 39528151
      9'hfe: T=64'b0111111111111101100010000101100100000001100100100001110100100000;  // 2147321945 26352928
      9'hff: T=64'b0111111111111111011000100001010100000000110010010000111110001000;  // 2147443221 13176712
      9'h100: T=64'b0111111111111111111111111111111100000000000000000000000000000000;  // 2147483647     0
      9'h101: T=64'b0111111111111111011000100001010111111111001101101111000001111000;  // 2147443221 -13176712
      9'h102: T=64'b0111111111111101100010000101100111111110011011011110001011100000;  // 2147321945 -26352928
      9'h103: T=64'b0111111111111010011100101101000011111101101001001101100100101001;  // 2147119824 -39528151
      9'h104: T=64'b0111111111110110001000011000000111111100110110111101010101000001;  // 2146836865 -52701887
      9'h105: T=64'b0111111111110000100101000111011111111100000100101101100100011010;  // 2146473079 -65873638
      9'h106: T=64'b0111111111101001110010111011111111111011010010011110011010100011;  // 2146028479 -79042909
      9'h107: T=64'b0111111111100001110001110110101011111010100000001111111111001011;  // 2145503082 -92209205
      9'h108: T=64'b0111111111011000100001111000110111111001101110000010011010000100;  // 2144896909 -105372028
      9'h109: T=64'b0111111111001110000011000011110111111000111011110101110010111011;  // 2144209981 -118530885
      9'h10a: T=64'b0111111111000010010101011001010111111000001001101010010001100010;  // 2143442325 -131685278
      9'h10b: T=64'b0111111110110101011000111011001011110111010111011111111101100110;  // 2142593970 -144834714
      9'h10c: T=64'b0111111110100111001101101011001111110110100101010110111110110111;  // 2141664947 -157978697
      9'h10d: T=64'b0111111110010111110011101011110011110101110011001111011101000100;  // 2140655292 -171116732
      9'h10e: T=64'b0111111110000111001010111111001011110101000001001001011111111011;  // 2139565042 -184248325
      9'h10f: T=64'b0111111101110101010011100111111111110100001111000101001111001011;  // 2138394239 -197372981
      9'h110: T=64'b0111111101100010001101101000111011110011011101000010110010100010;  // 2137142926 -210490206
      9'h111: T=64'b0111111101001101111001000101000011110010101011000010010001101110;  // 2135811152 -223599506
      9'h112: T=64'b0111111100111000010101111111010111110001111001000011110100011100;  // 2134398965 -236700388
      9'h113: T=64'b0111111100100001100100011011001111110001000111000111100010011010;  // 2132906419 -249792358
      9'h114: T=64'b0111111100001001100100011100001111110000010101001101100011010101;  // 2131333571 -262874923
      9'h115: T=64'b0111111011110000010110000101111111101111100011010101111110111000;  // 2129680479 -275947592
      9'h116: T=64'b0111111011010101111001011100010111101110110001100000111100110001;  // 2127947205 -289009871
      9'h117: T=64'b0111111010111010001110100011100011101101111111101110100100101011;  // 2126133816 -302061269
      9'h118: T=64'b0111111010011101010101011111101111101101001101111110111110010010;  // 2124240379 -315101294
      9'h119: T=64'b0111111001111111001110010101011011101100011100010010010001001111;  // 2122266966 -328129457
      9'h11a: T=64'b0111111001011111111001001001001011101011101010101000100101001111;  // 2120213650 -341145265
      9'h11b: T=64'b0111111000111111010101111111111011101010111001000010000001111011;  // 2118080510 -354148229
      9'h11c: T=64'b0111111000011101100100111110100111101010000111011110101110111100;  // 2115867625 -367137860
      9'h11d: T=64'b0111110111111010100110001010011111101001010101111110110011111011;  // 2113575079 -380113669
      9'h11e: T=64'b0111110111010110011001101000111011101000100100100010011000100010;  // 2111202958 -393075166
      9'h11f: T=64'b0111110110110000111111011111011111100111110011001001100100011000;  // 2108751351 -406021864
      9'h120: T=64'b0111110110001010010111110011111111100111000001110100011111000100;  // 2106220351 -418953276
      9'h121: T=64'b0111110101100010100010101100010111100110010000100011010000001101;  // 2103610053 -431868915
      9'h122: T=64'b0111110100111001100000001110101111100101011111010101111111011011;  // 2100920555 -444768293
      9'h123: T=64'b0111110100001111010000100001011111100100101110001100110100010001;  // 2098151959 -457650927
      9'h124: T=64'b0111110011100011110011101011000111100011111101000111110110010110;  // 2095304369 -470516330
      9'h125: T=64'b0111110010110111001001110010001111100011001100000111001101001101;  // 2092377891 -483364019
      9'h126: T=64'b0111110010001001010010111101110111100010011011001011000000011011;  // 2089372637 -496193509
      9'h127: T=64'b0111110001011010001111010100111111100001101010010011010111100010;  // 2086288719 -509004318
      9'h128: T=64'b0111110000101001111110111110110111100000111001100000011010000101;  // 2083126253 -521795963
      9'h129: T=64'b0111101111111000100010000010111111100000001000110010001111100101;  // 2079885359 -534567963
      9'h12a: T=64'b0111101111000101111000101000111111011111011000001000111111100100;  // 2076566159 -547319836
      9'h12b: T=64'b0111101110010010000010111000100011011110100111100100110001100001;  // 2073168776 -560051103
      9'h12c: T=64'b0111101101011101000000111001110111011101110111000101101100111011;  // 2069693341 -572761285
      9'h12d: T=64'b0111101100100110110010110100111011011101000110101011111001010001;  // 2066139982 -585449903
      9'h12e: T=64'b0111101011101111011000110010001111011100010110010111011110000010;  // 2062508835 -598116478
      9'h12f: T=64'b0111101010110110110010111010001111011011100110001000100010101001;  // 2058800035 -610760535
      9'h130: T=64'b0111101001111101000001010101101011011010110101111111001110100011;  // 2055013722 -623381597
      9'h131: T=64'b0111101001000010000100001101100011011010000101111011101001001010;  // 2051150040 -635979190
      9'h132: T=64'b0111101000000101111011101010110011011001010101111101111001111011;  // 2047209132 -648552837
      9'h133: T=64'b0111100111001000100111110110110111011000100110000110001000001100;  // 2043191149 -661102068
      9'h134: T=64'b0111100110001010001000111011000011010111110110010100011011011000;  // 2039096240 -673626408
      9'h135: T=64'b0111100101001010011111000001000111010111000110101000111010110110;  // 2034924561 -686125386
      9'h136: T=64'b0111100100001001101010010010110011010110010111000011101101111011;  // 2030676268 -698598533
      9'h137: T=64'b0111100011000111101010111010000111010101100111100100111011111111;  // 2026351521 -711045377
      9'h138: T=64'b0111100010000100100001000001001111010100111000001100101100010101;  // 2021950483 -723465451
      9'h139: T=64'b0111100001000000001100110010100011010100001000111011000110010001;  // 2017473320 -735858287
      9'h13a: T=64'b0111011111111010101110011000100011010011011001110000010001000110;  // 2012920200 -748223418
      9'h13b: T=64'b0111011110110100000101111101111111010010101010101100010100000101;  // 2008291295 -760560379
      9'h13c: T=64'b0111011101101100010011101101101011010001111011101111010110011110;  // 2003586778 -772868706
      9'h13d: T=64'b0111011100100011010111110010110011010001001100111001011111100010;  // 1998806828 -785147934
      9'h13e: T=64'b0111011011011001010010011000100011010000011110001010110110011110;  // 1993951624 -797397602
      9'h13f: T=64'b0111011010001110000011101010010111001111101111100011100010100000;  // 1989021349 -809617248
      9'h140: T=64'b0111011001000001101011110011110011001111000001000011101010110011;  // 1984016188 -821806413
      9'h141: T=64'b0111010111110100001011000000101011001110010010101011010110100011;  // 1978936330 -833964637
      9'h142: T=64'b0111010110100101100001011100111011001101100100011010101100111001;  // 1973781966 -846091463
      9'h143: T=64'b0111010101010101101111010100101111001100110110010001110100111110;  // 1968553291 -858186434
      9'h144: T=64'b0111010100000100110100110100010011001100001000010000110101111001;  // 1963250500 -870249095
      9'h145: T=64'b0111010010110010110010001000001111001011011010010111110110110001;  // 1957873795 -882278991
      9'h146: T=64'b0111010001011111100111011101000011001010101100100110111110101010;  // 1952423376 -894275670
      9'h147: T=64'b0111010000001011010100111111101011001001111110111110010100100111;  // 1946899450 -906238681
      9'h148: T=64'b0111001110110101111010111101000011001001010001011101111111101101;  // 1941302224 -918167571
      9'h149: T=64'b0111001101011111011001100010010111001000100100000110000110111010;  // 1935631909 -930061894
      9'h14a: T=64'b0111001100000111110000111100111111000111110110110110110001010000;  // 1929888719 -941921200
      9'h14b: T=64'b0111001010101111000001011010011011000111001001110000000101101101;  // 1924072870 -953745043
      9'h14c: T=64'b0111001001010101001011001000010011000110011100110010001011001110;  // 1918184580 -965532978
      9'h14d: T=64'b0111000111111010001110010100100011000101101111111101001000101111;  // 1912224072 -977284561
      9'h14e: T=64'b0111000110011110001011001101000111000101000011010001000101001001;  // 1906191569 -988999351
      9'h14f: T=64'b0111000101000001000010000000010011000100010110101110000111010111;  // 1900087300 -1000676905
      9'h150: T=64'b0111000011100010110010111100010111000011101010010100010110010000;  // 1893911493 -1012316784
      9'h151: T=64'b0111000010000011011110001111111011000010111110000011111000101011;  // 1887664382 -1023918549
      9'h152: T=64'b0111000000100011000100001001100111000010010001111100110101011011;  // 1881346201 -1035481765
      9'h153: T=64'b0110111111000001100100111000010011000001100101111111010011010100;  // 1874957188 -1047005996
      9'h154: T=64'b0110111101011111000000101011000111000000111010001011011001001001;  // 1868497585 -1058490807
      9'h155: T=64'b0110111011111011010111110001000111000000001110100001001101101001;  // 1861967633 -1069935767
      9'h156: T=64'b0110111010010110101010011001110010111111100011000000110111100011;  // 1855367580 -1081340445
      9'h157: T=64'b0110111000110000111000110100100110111110110111101010011101100110;  // 1848697673 -1092704410
      9'h158: T=64'b0110110111001010000011010001010010111110001100011110000110011100;  // 1841958164 -1104027236
      9'h159: T=64'b0110110101100010001001111111100110111101100001011011111000110000;  // 1835149305 -1115308496
      9'h15a: T=64'b0110110011111001001101001111101110111100110110100011111011001011;  // 1828271355 -1126547765
      9'h15b: T=64'b0110110010001111001101010001101110111100001011110110010100010100;  // 1821324571 -1137744620
      9'h15c: T=64'b0110110000100100001010010101111110111011100001010011001010110000;  // 1814309215 -1148898640
      9'h15d: T=64'b0110101110111000000100101101000010111010110110111010100101000100;  // 1807225552 -1160009404
      9'h15e: T=64'b0110101101001010111100100111100010111010001100101100101001110001;  // 1800073848 -1171076495
      9'h15f: T=64'b0110101011011100110010010110010010111001100010101001011111011001;  // 1792854372 -1182099495
      9'h160: T=64'b0110101001101101100110001010001110111000111000110001001100011010;  // 1785567395 -1193077990
      9'h161: T=64'b0110100111111101011000010100101010111000001111000011110111010010;  // 1778213194 -1204011566
      9'h162: T=64'b0110100110001100001001000110101110110111100101100001100110011100;  // 1770792043 -1214899812
      9'h163: T=64'b0110100100011001111000110001111110110110111100001010100000010010;  // 1763304223 -1225742318
      9'h164: T=64'b0110100010100110100111101000000010110110010010111110101011001101;  // 1755750016 -1236538675
      9'h165: T=64'b0110100000110010010101111010101010110101101001111110001101100011;  // 1748129706 -1247288477
      9'h166: T=64'b0110011110111101000011111011110010110101000001001001001101101001;  // 1740443580 -1257991319
      9'h167: T=64'b0110011101000110110001111101011110110100011000011111110001110001;  // 1732691927 -1268646799
      9'h168: T=64'b0110011011001111100000010001111110110011110000000010000000001101;  // 1724875039 -1279254515
      9'h169: T=64'b0110011001010111001111001011101110110011000111101111111111001100;  // 1716993211 -1289814068
      9'h16a: T=64'b0110010111011101111110111101001010110010011111101001110100111101;  // 1709046738 -1300325059
      9'h16b: T=64'b0110010101100011101111111001000110110001110111101111100111101001;  // 1701035921 -1310787095
      9'h16c: T=64'b0110010011101000100010010010010110110001010000000001011101011100;  // 1692961061 -1321199780
      9'h16d: T=64'b0110010001101100010110011011111110110000101000011111011100011110;  // 1684822463 -1331562722
      9'h16e: T=64'b0110001111101111001100101000111110110000000001001001101010110100;  // 1676620431 -1341875532
      9'h16f: T=64'b0110001101110001000101001100110010101111011010000000001110100010;  // 1668355276 -1352137822
      9'h170: T=64'b0110001011110010000000011010110010101110110011000011001101101100;  // 1660027308 -1362349204
      9'h171: T=64'b0110001001110001111110100110100010101110001100010010101110010010;  // 1651636840 -1372509294
      9'h172: T=64'b0110000111110001000000000011111010101101100101101110110110010010;  // 1643184190 -1382617710
      9'h173: T=64'b0110000101101111000101000110101110101100111111010111101011101001;  // 1634669675 -1392674071
      9'h174: T=64'b0110000011101100001110000010111110101100011001001101010100010001;  // 1626093615 -1402677999
      9'h175: T=64'b0110000001101000011011001100111010101011110011001111110110000011;  // 1617456334 -1412629117
      9'h176: T=64'b0101111111100011101100111000110110101011001101011111010110110110;  // 1608758157 -1422527050
      9'h177: T=64'b0101111101011110000011011011001010101010100111111011111100011110;  // 1599999410 -1432371426
      9'h178: T=64'b0101111011010111011111001000100110101010000010100101101100101110;  // 1591180425 -1442161874
      9'h179: T=64'b0101111001010000000000010101110110101001011101011100101101010111;  // 1582301533 -1451898025
      9'h17a: T=64'b0101110111000111100111010111101110101000111000100001000100000111;  // 1573363067 -1461579513
      9'h17b: T=64'b0101110100111110010100100011011010101000010011110010110110101011;  // 1564365366 -1471205973
      9'h17c: T=64'b0101110010110100001000001101111110100111101111010010001010101100;  // 1555308767 -1480777044
      9'h17d: T=64'b0101110000101001000010101100110010100111001010111111000101110100;  // 1546193612 -1490292364
      9'h17e: T=64'b0101101110011101000100010101001110100110100110111001101101101001;  // 1537020243 -1499751575
      9'h17f: T=64'b0101101100010000001101011100111010100110000011000010000111101110;  // 1527789006 -1509154322
      9'h180: T=64'b0101101010000010011110011001100110100101011111011000011001100111;  // 1518500249 -1518500249
      9'h181: T=64'b0101100111110011110111100001001010100100111011111100101000110010;  // 1509154322 -1527789006
      9'h182: T=64'b0101100101100100011001001001011110100100011000101110111010101101;  // 1499751575 -1537020243
      9'h183: T=64'b0101100011010100000011101000110010100011110101101111010100110100;  // 1490292364 -1546193612
      9'h184: T=64'b0101100001000010110111010101010010100011010010111101111100100001;  // 1480777044 -1555308767
      9'h185: T=64'b0101011110110000110100100101010110100010110000011010110111001010;  // 1471205973 -1564365366
      9'h186: T=64'b0101011100011101111011101111100110100010001110000110001010000101;  // 1461579513 -1573363067
      9'h187: T=64'b0101011010001010001101001010100110100001101011111111111010100011;  // 1451898025 -1582301533
      9'h188: T=64'b0101010111110101101001001101001010100001001010001000001101110111;  // 1442161874 -1591180425
      9'h189: T=64'b0101010101100000010000001110001010100000101000011111001001001110;  // 1432371426 -1599999410
      9'h18a: T=64'b0101010011001010000010100100101010100000000111000100110001110011;  // 1422527050 -1608758157
      9'h18b: T=64'b0101010000110011000000100111110110011111100101111001001100110010;  // 1412629117 -1617456334
      9'h18c: T=64'b0101001110011011001010101110111110011111000100111100011111010001;  // 1402677999 -1626093615
      9'h18d: T=64'b0101001100000010100001010001011110011110100100001110101110010101;  // 1392674071 -1634669675
      9'h18e: T=64'b0101001001101001000100100110111010011110000011101111111111000010;  // 1382617710 -1643184190
      9'h18f: T=64'b0101000111001110110101000110111010011101100011100000010110011000;  // 1372509294 -1651636840
      9'h190: T=64'b0101000100110011110011001001010010011101000011011111111001010100;  // 1362349204 -1660027308
      9'h191: T=64'b0101000010010111111111000101111010011100100011101110101100110100;  // 1352137822 -1668355276
      9'h192: T=64'b0100111111111011011001010100110010011100000100001100110101110001;  // 1341875532 -1676620431
      9'h193: T=64'b0100111101011110000010001110001010011011100100111010011001000001;  // 1331562722 -1684822463
      9'h194: T=64'b0100111010111111111010001010010010011011000101110111011011011011;  // 1321199780 -1692961061
      9'h195: T=64'b0100111000100001000001100001011110011010100111000100000001101111;  // 1310787095 -1701035921
      9'h196: T=64'b0100110110000001011000101100001110011010001000100000010000101110;  // 1300325059 -1709046738
      9'h197: T=64'b0100110011100001000000000011010010011001101010001100001101000101;  // 1289814068 -1716993211
      9'h198: T=64'b0100110000111111110111111111001110011001001100000111111011100001;  // 1279254515 -1724875039
      9'h199: T=64'b0100101110011110000000111000111110011000101110010011100000101001;  // 1268646799 -1732691927
      9'h19a: T=64'b0100101011111011011011001001011110011000010000101111000001000100;  // 1257991319 -1740443580
      9'h19b: T=64'b0100101001011000000111001001110110010111110011011010100001010110;  // 1247288477 -1748129706
      9'h19c: T=64'b0100100110110100000101010011001110010111010110010110000110000000;  // 1236538675 -1755750016
      9'h19d: T=64'b0100100100001111010101111110111010010110111001100001110011100001;  // 1225742318 -1763304223
      9'h19e: T=64'b0100100001101001111001100110010010010110011100111101101110010101;  // 1214899812 -1770792043
      9'h19f: T=64'b0100011111000011110000100010111010010110000000101001111010110110;  // 1204011566 -1778213194
      9'h1a0: T=64'b0100011100011100111011001110011010010101100100100110011101011101;  // 1193077990 -1785567395
      9'h1a1: T=64'b0100011001110101011010000010011110010101001000110011011010011100;  // 1182099495 -1792854372
      9'h1a2: T=64'b0100010111001101001101011000111110010100101101010000110110001000;  // 1171076495 -1800073848
      9'h1a3: T=64'b0100010100100100010101101011110010010100010001111110110100110000;  // 1160009404 -1807225552
      9'h1a4: T=64'b0100010001111010110011010101000010010011110110111101011010100001;  // 1148898640 -1814309215
      9'h1a5: T=64'b0100001111010000100110101110110010010011011100001100101011100101;  // 1137744620 -1821324571
      9'h1a6: T=64'b0100001100100101110000010011010110010011000001101100101100000101;  // 1126547765 -1828271355
      9'h1a7: T=64'b0100001001111010010000011101000010010010100111011101100000000111;  // 1115308496 -1835149305
      9'h1a8: T=64'b0100000111001110000111100110010010010010001101011111001011101100;  // 1104027236 -1841958164
      9'h1a9: T=64'b0100000100100001010110001001101010010001110011110001110010110111;  // 1092704410 -1848697673
      9'h1aa: T=64'b0100000001110011111100100001110110010001011010010101011001100100;  // 1081340445 -1855367580
      9'h1ab: T=64'b0011111111000101111011001001011110010001000001001010000011101111;  // 1069935767 -1861967633
      9'h1ac: T=64'b0011111100010111010010011011011110010000101000001111110101001111;  // 1058490807 -1868497585
      9'h1ad: T=64'b0011111001101000000010110010110010010000001111100110110001111100;  // 1047005996 -1874957188
      9'h1ae: T=64'b0011110110111000001100101010010110001111110111001110111101100111;  // 1035481765 -1881346201
      9'h1af: T=64'b0011110100000111110000011101010110001111011111001000011100000010;  // 1023918549 -1887664382
      9'h1b0: T=64'b0011110001010110101110100111000010001111000111010011010000111011;  // 1012316784 -1893911493
      9'h1b1: T=64'b0011101110100101000111100010100110001110101111101111011111111100;  // 1000676905 -1900087300
      9'h1b2: T=64'b0011101011110010111011101011011110001110011000011101001100101111;  // 988999351 -1906191569
      9'h1b3: T=64'b0011101001000000001011011101000110001110000001011100011010111000;  // 977284561 -1912224072
      9'h1b4: T=64'b0011100110001100110111010011001010001101101010101101001101111100;  // 965532978 -1918184580
      9'h1b5: T=64'b0011100011011000111111101001001110001101010100001111101001011010;  // 953745043 -1924072870
      9'h1b6: T=64'b0011100000100100100100111011000010001100111110000011110000110001;  // 941921200 -1929888719
      9'h1b7: T=64'b0011011101101111100111100100011010001100101000001001100111011011;  // 930061894 -1935631909
      9'h1b8: T=64'b0011011010111010001000000001001110001100010010100001010000110000;  // 918167571 -1941302224
      9'h1b9: T=64'b0011011000000100000110101101100110001011111101001010110000000110;  // 906238681 -1946899450
      9'h1ba: T=64'b0011010101001101100100000101011010001011101000000110001000110000;  // 894275670 -1952423376
      9'h1bb: T=64'b0011010010010110100000100100111110001011010011010011011101111101;  // 882278991 -1957873795
      9'h1bc: T=64'b0011001111011110111100101000011110001010111110110010110010111100;  // 870249095 -1963250500
      9'h1bd: T=64'b0011001100100110111000101100001010001010101010100100001010110101;  // 858186434 -1968553291
      9'h1be: T=64'b0011001001101110010101001100011110001010010110100111101000110010;  // 846091463 -1973781966
      9'h1bf: T=64'b0011000110110101010010100101110110001010000010111101001111110110;  // 833964637 -1978936330
      9'h1c0: T=64'b0011000011111011110001010100110110001001101111100101000011000100;  // 821806413 -1984016188
      9'h1c1: T=64'b0011000001000001110001110110000010001001011100011111000101011011;  // 809617248 -1989021349
      9'h1c2: T=64'b0010111110000111010100100110001010001001001001101011011001111000;  // 797397602 -1993951624
      9'h1c3: T=64'b0010111011001100011010000001111010001000110111001010000011010100;  // 785147934 -1998806828
      9'h1c4: T=64'b0010111000010001000010100110001010001000100100111011000100100110;  // 772868706 -2003586778
      9'h1c5: T=64'b0010110101010101001110101111101110001000010010111110100000100001;  // 760560379 -2008291295
      9'h1c6: T=64'b0010110010011000111110111011101010001000000001010100011001111000;  // 748223418 -2012920200
      9'h1c7: T=64'b0010101111011100010011100110111110000111101111111100110011011000;  // 735858287 -2017473320
      9'h1c8: T=64'b0010101100011111001101001110101110000111011110110111101111101101;  // 723465451 -2021950483
      9'h1c9: T=64'b0010101001100001101100010000000110000111001110000101010001011111;  // 711045377 -2026351521
      9'h1ca: T=64'b0010100110100011110001001000010110000110111101100101011011010100;  // 698598533 -2030676268
      9'h1cb: T=64'b0010100011100101011100010100101010000110101101011000001111101111;  // 686125386 -2034924561
      9'h1cc: T=64'b0010100000100110101110010010100010000110011101011101110001010000;  // 673626408 -2039096240
      9'h1cd: T=64'b0010011101100111100111011111010010000110001101110110000010010011;  // 661102068 -2043191149
      9'h1ce: T=64'b0010011010101000001000011000010110000101111110100001000101010100;  // 648552837 -2047209132
      9'h1cf: T=64'b0010010111101000010001011011011010000101101111011110111100101000;  // 635979190 -2051150040
      9'h1d0: T=64'b0010010100101000000011000101110110000101100000101111101010100110;  // 623381597 -2055013722
      9'h1d1: T=64'b0010010001100111011101110101011110000101010010010011010001011101;  // 610760535 -2058800035
      9'h1d2: T=64'b0010001110100110100010000111111010000101000100001001110011011101;  // 598116478 -2062508835
      9'h1d3: T=64'b0010001011100101010000011010111110000100110110010011010010110010;  // 585449903 -2066139982
      9'h1d4: T=64'b0010001000100011101001001100010110000100101000101111110001100011;  // 572761285 -2069693341
      9'h1d5: T=64'b0010000101100001101100111001111110000100011011011111010001111000;  // 560051103 -2073168776
      9'h1d6: T=64'b0010000010011111011100000001110010000100001110100001110101110001;  // 547319836 -2076566159
      9'h1d7: T=64'b0001111111011100110111000001101110000100000001110111011111010001;  // 534567963 -2079885359
      9'h1d8: T=64'b0001111100011001111110010111101110000011110101100000010000010011;  // 521795963 -2083126253
      9'h1d9: T=64'b0001111001010110110010100001111010000011101001011100001010110001;  // 509004318 -2086288719
      9'h1da: T=64'b0001110110010011010011111110010110000011011101101011010000100011;  // 496193509 -2089372637
      9'h1db: T=64'b0001110011001111100011001011001110000011010010001101100011011101;  // 483364019 -2092377891
      9'h1dc: T=64'b0001110000001011100000100110101010000011000111000011000101001111;  // 470516330 -2095304369
      9'h1dd: T=64'b0001101101000111001100101110111110000010111100001011110111101001;  // 457650927 -2098151959
      9'h1de: T=64'b0001101010000010101000000010010110000010110001100111111100010101;  // 444768293 -2100920555
      9'h1df: T=64'b0001100110111101110010111111001110000010100111010111010100111011;  // 431868915 -2103610053
      9'h1e0: T=64'b0001100011111000101110000011110010000010011101011010000011000001;  // 418953276 -2106220351
      9'h1e1: T=64'b0001100000110011011001101110100010000010010011110000001000001001;  // 406021864 -2108751351
      9'h1e2: T=64'b0001011101101101110110011101111010000010001010011001100101110010;  // 393075166 -2111202958
      9'h1e3: T=64'b0001011010101000000100110000010110000010000001010110011101011001;  // 380113669 -2113575079
      9'h1e4: T=64'b0001010111100010000101000100010010000001111000100110110000010111;  // 367137860 -2115867625
      9'h1e5: T=64'b0001010100011011110111111000010110000001110000001010100000000010;  // 354148229 -2118080510
      9'h1e6: T=64'b0001010001010101011101101011000110000001101000000001101101101110;  // 341145265 -2120213650
      9'h1e7: T=64'b0001001110001110110110111011000110000001100000001100011010101010;  // 328129457 -2122266966
      9'h1e8: T=64'b0001001011001000000100000110111010000001011000101010101000000101;  // 315101294 -2124240379
      9'h1e9: T=64'b0001001000000001000101101101010110000001010001011100010111001000;  // 302061269 -2126133816
      9'h1ea: T=64'b0001000100111001111100001100111110000001001010100001101000111011;  // 289009871 -2127947205
      9'h1eb: T=64'b0001000001110010101000000100100010000001000011111010011110100001;  // 275947592 -2129680479
      9'h1ec: T=64'b0000111110101011001001110010101110000000111101100110111000111101;  // 262874923 -2131333571
      9'h1ed: T=64'b0000111011100011100001110110011010000000110111100110111001001101;  // 249792358 -2132906419
      9'h1ee: T=64'b0000111000011011110000101110010010000000110001111010100000001011;  // 236700388 -2134398965
      9'h1ef: T=64'b0000110101010011110110111001001010000000101100100001101110110000;  // 223599506 -2135811152
      9'h1f0: T=64'b0000110010001011110100110101111010000000100111011100100101110010;  // 210490206 -2137142926
      9'h1f1: T=64'b0000101111000011101011000011010110000000100010101011000110000001;  // 197372981 -2138394239
      9'h1f2: T=64'b0000101011111011011010000000010110000000011110001101010000001110;  // 184248325 -2139565042
      9'h1f3: T=64'b0000101000110011000010001011110010000000011010000011000101000100;  // 171116732 -2140655292
      9'h1f4: T=64'b0000100101101010100100000100100110000000010110001100100101001101;  // 157978697 -2141664947
      9'h1f5: T=64'b0000100010100010000000001001101010000000010010101001110001001110;  // 144834714 -2142593970
      9'h1f6: T=64'b0000011111011001010110111001111010000000001111011010101001101011;  // 131685278 -2143442325
      9'h1f7: T=64'b0000011100010000101000110100010110000000001100011111001111000011;  // 118530885 -2144209981
      9'h1f8: T=64'b0000011001000111110110010111110010000000001001110111100001110011;  // 105372028 -2144896909
      9'h1f9: T=64'b0000010101111111000000000011010110000000000111100011100010010110;  // 92209205 -2145503082
      9'h1fa: T=64'b0000010010110110000110010101110110000000000101100011010001000001;  // 79042909 -2146028479
      9'h1fb: T=64'b0000001111101101001001101110011010000000000011110110101110001001;  // 65873638 -2146473079
      9'h1fc: T=64'b0000001100100100001010101011111110000000000010011101111001111111;  // 52701887 -2146836865
      9'h1fd: T=64'b0000001001011011001001101101011110000000000001011000110100110000;  // 39528151 -2147119824
      9'h1fe: T=64'b0000000110010010000111010010000010000000000000100111011110100111;  // 26352928 -2147321945
      9'h1ff: T=64'b0000000011001001000011111000100010000000000000001001110111101011;  // 13176712 -2147443221
      default: T=64'b0;
    endcase

endmodule
